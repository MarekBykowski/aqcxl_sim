`protected

    MTI!#?GYx1Dx#O!wnvKe'j]_Tc];G\xz_R\o3[Q3\w|.,.}3r-^I#s!YxG!]+uB\'Xk5W]<[QZk{
    MaDTZl511VZ^i%13C~E*ve!{lQ[C~~;>e?=V_^$_$1jIxEIRG_=BKZq?XXvVz<Q.pL$?~7A-e#>T
    ]z}Uz$2R,KkR!n$wT5l*n~Z]Hn>{AE2awlQa;l{,'*Msx,Ew]v!QGi{SF&m-+{p=*KND~DrweK?h
`endprotected
