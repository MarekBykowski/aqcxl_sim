`protected

    MTI!#*Y^IWX![\!z#~GlGOAB{0];G\xz_R\rn[Q3\w|.[rXjj5z=Yjj#Jjm*<aAj'><CeivT>}r"
    qwE-Z>a,jY^?Rw=]-1}~?^H-_BnoRin;e0L=~aInEZ,5Ky>7-2'Cn>2I'atm5vQ_HAexz^@oG[zB
    ''Q77@Gt{V>$Pil|.Cn3$I5!o|%j-BA-eAn7?ju;r7#{Ek]yN,e\ndX=?nW-uj=#2]V3l17+UEa{
    dZTXkFIET$NkvDrQV^kB517ir1BQ[1-envp!|npm>'V+kHD-z=bw5Yw=XA3EG!W\3xW|\WDBk{!^
    Y}?_]$_rz}Hwa<j!%[mCls<TKRGVYk-E}[uZD]OWHDHJ@D3'R=HxR$<+Gk}}-><BC+jm-@[i_51Q
    1$C!Q=@[Rjl?HX5$BH+3^|{[mOx*-Br][;DaDBKOr+C_s'{<l?-]'[Qz'CfeA=p7sz=8Y#\z={]\
    7:PW'jQE~{vZCXZs$p!=\BJ9[eZA=E*}C5eO_7j;/]_[i__7+7Z{K!H!jWRU[c9'EeKeOT
`endprotected
