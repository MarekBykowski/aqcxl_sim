`protect
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_2)
//pragma protect key_method=RSA
//pragma protect key_block
AOo66z1Sgv/a9QvgH5q3RKtkumNo4YfjdnPEgyHg8uc/M2G+JRIbSeRbubj3sDn3
STVBTVxFAHptkaNCdotBqX/NULh7JQow0MLNUBsgKduC3tb2PI931copwIma8YcR
g8+no3G5l63lfEiS7SA0YlHKhHOsEivd2mFeBSQnTGHDhpzifpC9GKx1WTgS4tea
R4rs9mex0HoIuyWRjhYyTi+YqmBvNqelFYGjcFD1+/AvNJ6LDW+kGalMycQ19LaT
SDdXHZN+kwvycH5/FSWyQqzzxf/Zl3mNooQ7ZO9xi3myNstxJ4P1lvwhfnlg1e5I
ozmKNCPGQP3P37A2T4Kshg==
//pragma protect end_key_block
//pragma protect digest_block
MtcXbWjW3EKUtHpGuKvF4r8B+iU=
//pragma protect end_digest_block
//pragma protect data_block
H0HJd7wFB5Fv86WT6dj9Ju/sKMhvpRFnFTySenwfwGaUp6/FXWDcE4qLe/vsDdIy
qeQo/fGH8M0pCxs5tQ7+saO3AUKX6Ar0pr7DF9fGu1zs4dBgeiB76RClMfdlcD+n
NkQ2X9kxAHxuqKoolocfbbWnLpPpPdzMPhTfJP5MpuQV+hth3A/obv7jB4sbAi+6
CMb5GKbNVhwvWtmaez2+xLfzayGTBmKica79OeRVEwk4qOVJpUWAUXSJyZgkIzM4
3wM2TkhV0gnopxkaVvYYZ1+lWSqfwU/nSpedQwG4rmi8U12TyjIkrUfcVqGxeFiN
ODub2YazrL3bIwVZm1T4j2sF4sBJGw+Agx5004U5QEO7PZDWwkBYvisBmJX2JtJG
r6p1RTeSLrzu08FKaMjG8FQDHkcr7o2htXr419csyxijWhZ1/JJ4fapxJF4HPoyN
//pragma protect end_data_block
//pragma protect digest_block
ykQQKWZTw5UcJjhPsCtSaYcPRGY=
//pragma protect end_digest_block
//pragma protect end_protected
    `include "qemu_enum.svh"
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_2)
//pragma protect key_method=RSA
//pragma protect key_block
Aly9ogwPRyDI8/iZGAEOSu4n15rK6UfhCxyaX+6PqsliJBdzShteUjqm8RZop7Xd
cI0GvXmW9Zyr7DxMnTB8lRC79bKyOpkhRujME/dKJ1dC94flpmpQpoQNMy5MeqtJ
JgWWPICyMN5L5ydvDHuSmsKVbHFVVTMj6R7lq+P66MZYguppjAB2vCJIuto1vw0c
1UkIDSefeYUTmOOLjTwo9YpWNlAV3I4V9Sz3FjuB1Pzx4R5cUQsYpL11edqLLLcO
Z+6YCFYQi0zZrMsSA61Z8n3jTYhVVoPEGe8sm9Txriy9es6bvGvPrR0BqJfSn3E5
0wWQYvyfok/cM7bgzuCc4g==
//pragma protect end_key_block
//pragma protect digest_block
hkAZrYK4Td1imLpELfOKDVyUkJc=
//pragma protect end_digest_block
//pragma protect data_block
4Xu0hh6/x5Th3Y5U7m/iXuut8uvfxgxWbSQsb58btdMh8xzlfDlTbyeK8E2Dg0MS
ZfkWV8WTwBdNJuI8vYdm/gjEMP9lUkQTQ39Wopn5L/VWQXklbslbU2SxsEG1hsBx
C/EUasKPXXjmczYzZKdUO//6Iqz1QUa/Kc4ZCs8VCfl8pep2FkwixizRO0EuvSBi
Kx+7lbVXLlR8a8WG/FWKi4MAz+QSD2s+n4FkCX9+9KmE1+TemEgpfoa/ANRzYhO7
o6xhPhfIfSfD4vQjo1MfKPE87o1t1cCzzSrrXLUMnyrqH0ofGSatxmb0k6a5jjWt
t/aiIFPZEEmqItOY9Gwwv/HK1ny0vphL53oKtBu9wkEartRsAFlfezs00dJA8lTy
4Vgk7nGxMr1nqxiEx5pFHrOLm+BCiQCOL9fYi33epNJXVIipxgZu5WO3bO8R3mWk
3BBP4KLuBKTQmInWSIy3g1/DVcm+crVfFy42XAgIRwCiSQjprEClMDUatZJSWM6V
mdQ8qDCe6jP1T+ePO88Ozl2ILz+aVIzkcd/TvgXkYIjZnJo6pW0QYF9WgClXQCp0
B2VA7G9f4RJ7eXYub0pETtFyYFTZWhCifF2CcvOXIDnfbGxtjp3zrRZjy3wLe7BH
VbXjv0Xa5gPCCzm61u/oUY5ABmLKR42t23frAMA0Z/4rW6/xySFU/a9M1pYxSom7
wm7vT3MQELmoUXmr023BWwbrVot/drCgxImw8D2tlZTwP1Yc+pq+swam7KrgolcC
2qsz/bbo93gvmvQhgUx8JHDgChk1EXriNHm4iQsAznUGEG713IY66r2rL+7aTQn7
GTOc7hzvffyUseAJf94CjZZNZGvIOZSE5CgtYDUMiccoZwbiVjzyr5F6D46fnVi8
C2C0hkW8BqcbrU3CKOSqcxWVdnmTsIlC3x0gaG6cMAxoJwY0S9QMNfkTu/PZqu9b
32doyBeN4zhbgfDyXRxHuA==
//pragma protect end_data_block
//pragma protect digest_block
A4/N7Nrtn/xHQ0CkMsOFm8XClNo=
//pragma protect end_digest_block
//pragma protect end_protected
