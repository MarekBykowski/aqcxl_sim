package qemu_rx_pkg;
import avery_pkg::*;
import apci_pkg::*;
import apci_pkg_test::*;
import qemu_simc_pkg::*;

`include "qemu_enum.svh"
`ifdef INTEL_IOSF
`include "qemu_iosf.svh"
`endif
`ifdef AVERY_SPDM
`include "spdm_dpi.svh"
`endif
`include "measure.svh"

bit RST_TYPE = 0; // 1 for Hot 0 for Warm/Cold reset
bit PM_SUP = 0; // 1 for Power Management support
typedef bit[31:0] payload_t[$];
typedef apci_tlp acpi_tlp_q_t[$];
typedef payload_t addr_payload_hash_t[bit [63:0]];
typedef acpi_tlp_q_t addr_dropped_cpld_hash_t[bit [63:0]];
// size in bytes of the simcluster buffer
bit [31:0] qemu_debug_g= 3;
bit [31:0] vip_type_g= 0;
bit edb_logerror_jump_g= 0;
apci_tlp dropped_cpld_q[$];
addr_dropped_cpld_hash_t mrd_dropped_cpld_tlp;
addr_payload_hash_t mrd_dropped_cpld_payload;
bit[63 :0]  _all_one_64 = '1;
bit[63 :0]  _all_zero_64 = '0;
apci_atc_mgr atc_mgr;
bit[63:0] ats_xaddr;
bit[127:0] base_limit_Q[$];
bit[3:0] evict_mode = 4'b0011;
bit[63:0] max_clines = 8;
bit[11:0] pm_cap;
bit[11:0] exp_cap;
// Do not refactor PERST_N this is for sideband
bit PERST_N = 1; // active low
apci_device ep0;
apci_device all_bfms[$];
// use integer instead of int to avoid vpi issue
static integer aqemu_int1, aqemu_int3;

string sc_key= append_key_after_user(`simcluster_QEMU_key);
string edb_key= append_key_after_user(`simcluster_EDB_key);
`define SUBCMD_SHIFT (8)
`define CMD_MASK (8'hf)

`ifndef APCI_MPORT
`define PORT_NUM 1
`else
`define PORT_NUM 2
`endif

task automatic set_hdm_range(ref apci_device bfm);
    apci_bdf_t        hdm_bdf[`PORT_NUM];
    apci_addr_range_t hdm_ranges[`PORT_NUM][$];
    bit[63:0] ig = (1 << (8 + 6)); // 6 : 16 KB
    bit[63:0] iw = `PORT_NUM;
    bit[63:0] hdm_base = 64'h1_9000_0000;
    bit[63:0] hdm_len = 64'h0_4000_0000;

`ifdef AVERY_CXL_1_1
    hdm_bdf[0]  = 'h000;
`else
    for (int i = 0; i < `PORT_NUM; i++)
        hdm_bdf[i]  = (i + 1) * 'h100;
`endif

    /* Create RC HDM bkdoor mapping for single, 
     1 decoder 2 ep +APCI_MPORT
     2 decoder 2 ep +APCI_MPORT +SEPARATE_EP */
    if (`PORT_NUM == 1) begin
        apci_addr_range_t range;
        range.base = 64'h1_9000_0000;
        range.len =  64'h2000_0000;
        hdm_ranges[0].push_back(range);
    	bfm.cxl_bkdoor_add_hdm(0, hdm_ranges[0], hdm_bdf[0]);
    end
`ifdef SEPARATE_EP
    // for separate devices
    for (longint i = 0; i < `PORT_NUM; i++) begin
        apci_addr_range_t range;
        range.base = 64'h1_9000_0000 + 'h2000_0000 * i;
        range.len =  64'h2000_0000;
        hdm_ranges[i].push_back(range);
    end

    for (longint i = 0; i < `PORT_NUM; i++) begin
    	bfm.cxl_bkdoor_add_hdm(i, hdm_ranges[i], hdm_bdf[i]);
    end
`else
`ifdef APCI_MPORT
    // For iw == 2
    for (longint i = 0; i < (hdm_len / ig); i++) begin
        apci_addr_range_t range;
        range.base = hdm_base + i * ig;
        range.len = ig;
        hdm_ranges[(i % iw)].push_back(range);
    end
    for (int i = 0; i < `PORT_NUM; i++)
        bfm.cxl_bkdoor_add_hdm(i % iw, hdm_ranges[(i % iw)], hdm_bdf[(i % iw)]);
`endif // APCI_MPORT
`endif // SEPARATE_EP
endtask

`protected
L?;\WcAGEK^TQ&bULe-/=4ON\^/<3@:.P),g@LIff0=2f5NE/EF?()P\U1LaI7YG
^F2:A)[4N#gAJM-WN@-/E<FFaO)>;J/=D&J;bW@&3;/KJ?/01-)d<NX4<UbdXOQV
g<fU.1&<N0RKOGYAV;()LA#XCXDSHO#:<a)T(a^EX5(=@UWeK[V-S+&,=bONLBgI
cZ49gHASOEH,839\WFDJTB^-:9&,=83J.VaP[#cB=;QUOSW@.T_?gT@gFcQFM55/
,.CI7^1J+NK_F<-U-G<=;#GHbO1N)GV)3e3X(+[3;9L2bZ@M23ST:^<eS_\F-48+
U,C/;e[,\Gg66V]&=WGQP;1C?0Zg7Q^TEFE\SC[Y@eDFMa].>HIUMS\>5Bbf.<B=
-2XU99M8>@GMW0N#O=MA6dH<9W+Ia9L-U3J8&<2[.)2:K9<Fa(2Ad)WcPF:(40,H
;Hc^=5TLQRF\g=(ZD#J#3^)@JLN<?AQGBMeSgO35.U-ORZ9eEdB);J4UYY4IKcbW
AL78SQa5SNRbV324.+Mc)\/Sd0N92SNR.>PFRTPgIf_[=)V/FP,TW^WWN=_,<7Y)
5AG#1-F&HfLb(<a_=/-@-NXYTVKEAV[;e.cM9QcS+L.G3,9.TQ&50gKMU7f=;7K:
CW;Y[U#b].fYgH\fW5A&KY)]beGb&^CK#VW/bXCY97;CK&WTPbBI,Z2W,)f58:]c
d&Qa(K)0E:08A.4NH<;&UX8;b2Q^AUeUXga@+UJBg?9932@6XEA>F4TM.-T?-#K1
2?G5/]@Y4_3@c/=Bgd4O(9P9,V=.(&Z-MA0@^Na>e#M#)/GF)P=J97_:cb)f^[^A
J=\Da_.@>D)=/[KV_Rc]_M\C1VH<UN2^f[_eC\^_4QJ3gCT:7<bQM0(YU=6b+dLf
Pa0X/89^gd.MH2A;A@6b,\FG:OY]P_cJP=Jcgb<888a3F-N(Z:Ac/aAB>a(1b:V^
+E\a6Y7B?,]YMH<a&Keb8G(,OGZMDL-)OK\:8gH(;ORQ:\/0:b:B@6e^));C<U2e
1Eg/]@E.Pd>UG7Y1=_PeDTRSQIRb,R<0Dg2W9:;_\H5/>I](gT&5TD#PAC>^;=PK
;S3c?Ce;\LYAH/;W\\<SdHe/&45a()NSM83(-39TCVX;6.)K:ZgK_S4,G5?M#Db-
4S\JIcEV:cLAY,UH\F+:X-^aIa@PSdGX0&E2R+)+ZW58BWG_5:/Y]dA9B&13IS++
+1ZZEa&0Ka=D_N0D;2(Xb.7F?GIZ,JJ/@-eL4-R^+O,-.&_KZaH>\JYF1)4gL8E\
H)NNVHAIKb<^RdW.;VgFaK:D[#gd:C3C+;d\]=eKgV&_1gSVQP8)C549GW-0S3JL
V#9d75dP(D])])(f-8&+fcLM&BaZ>T]3BVO^\@D&.\cB,RfP[].L#E/d4X,?JfKX
6\MB1;[DJOe2:13C12(E7c:^5^\e/J0TBgPc5?0./bU6LY)ZPOU&=g2PQ0UOX7dQ
70b5?]24&H#]cY381Y1-HV<8c[_9FL^U42=b8A\ccaNS^)0AgQ6\7GOKTI/I\_/\
GM+7U?ZMO^b;XOSCMS@,9DLE>3\]W,WL)>D?@HT;RDGSbK;5I]^UB1)bgV:FUDLf
92NIA^d_Z:4[[O+<9GY6)\9E^Z-V24GcTP?^RE0D_GAO_&+O0_UNGSSCFADcB>=3
ZdQQ17PfONGAaPX4R060XJ?7AVXK,SU^4IF1Pe[^G[.M3G<6ObWc=.YfaL.JXUO?
YP^]^1;Q_35\0bZ//Cg[QOGgNLF,&;0P&;&K/6X7_KIgO#D\Sa(1(Z&XT+9@5M6(
((E9II?D6a&<Hf]X3A,T.N/GB^-&YdSOc;d/?]:9V)^_<7PR&e+Q(aMdb#N&#7a2
F2^bN3f#DEZF:)-1V>KZ9&N^Naa>E\[GIcP?V)g+Lb]WU0c>^+@Y^Q6XRed__UU0
Z-?B.7D)LRE03X>cYH&0^MH9.aBYGTgJ8a\XAZ+[Nb^#XWSF^7&J;FUQRQ/FUKGE
;4U.(RL#&#N)9>[BaMaTG-:T?&U_>Nb[GG+>>L22PLYcLUE6-X:cJ7d>F,Lc;Nc]
6\=\)&Q>7;\I7DcN/VX9F,896a#UFR=2>+A_9d]R8dMbA917LVD5Z;1#A2E@ZLBP
[E3?OKWE7&1=TQJT\0>XV+ZTHU:@c45VKJG]\9HML)G:;b23F5<7IRN)7<=N;Z)B
Z(4@PB1K>6_321YF>>ZPg\Ff_YX9,>_QFCZ>2PeCIBYU?W-5bf#X.:,/<:3C3YET
d@f2\NeQO+P?M&7;R<a#e-A8[I&9U3;3G1B-P^[BW,U]DfO5,_]J&1gDOO\^^YT6
(&B\K,^b[PPNK\GBX+>#_SPG4=E9(-.RF;HM;N-@QYMO2DPUY^X^(Z]:=ZM/;^7^
@@^B(ESF\9]P/KX/Mg5+TFT?0b4D?@J5)9Pg1[bUa7gdC89NdY4HS#F_747Y+ZU3
R[E(#_:b.3J5Q0VgESQIBC)=ObVa5.V=(?(Q+GX9g/5TD[F@0AHOS-cW7?YOd.E.
2X:\>L0OJYBON1R1ZF[_8)20)N)Q=L<a3dL5HT^1H)0QBT.(?,5;YQ>c-5bJ&\&4
\[OT7fG<R43Jd&EI?+aRXP2MJ4PF1Bg:EO=Q+]-;8]YWC_BJ);02XU5>FY0U?E,,
8B[4(e:-7L^NYU_>&I6F]C>.5C9D;LPe&e_E]TWRKU#0#V,+>LWKT,3O<,GL0XRX
C<^Yc7)?<EUc>@G5Q]E=Uf2Mb<GGU/@VWMPN,A,(Da8:a=>^L3D1^7Y-a&0T;</(
<TX981.,5dee#D5YaE-d0C4EK;,U9#QMSg/&MEJFS@Bg_d?-V31=\;E\:65@f@<Y
5ZGSO.QM<Y-dY72.,@<=H8Y&RW0S+/YQK@,eQ<N7\C(B(LPG=R.(g#\>O4,852Td
BA-HK0MIKP_1I<fEKU>e--)A)bQK1\KPX6(@2\E8X3/CHY.;b[)TA#cO]KR-MUDB
#@&K;DAP;_#DV-X)fA;Q.FL<OE#dffFO?ZZU:YSC^cJDcVUFc6P\Z:A]d1J(_718
aFKH3>4a)^f7\:c()@M8_<&?a1WKY0@c1GeaU7D-ZC42/N:A/FJ,EO.ZO&RDUI6:
#]e[f@GdPH6d:E5;S=3)g0&:Og6B:N(.d8TGXZ+_-.(1ST?H(5_OECI#<=BaO=42
&5POKPcOUCG/FS:FGHdD-&PY&7/OZVEFf3_C]?;PJVc_,+[J=X3:Z@gM<(EDK8Y^
_C<bT(8YUE(a_C@(N8GJCQYP)>?)-KBDfZ\<IJ4Q_g\b]J5?Q@f\T3.fN&?Og6-^
TbRVCeG72()1PYafKA_-76SE[fHQ#1+=3&9b[YV&(_FB[(Zdac.A:c&AL0)>W6<?
KF5?;:@)UMHFSd;Oc)[SMND,0+(R0BRHcYf5a]D1B&;9;SSQ>cIMc]P^9G4bVBfJ
BPX[)TZ_Y#/57FR2,+?)E-aJ]/S\MS28X>CU+S>GcV-O\\/=?#fS>NHcJ\+>#[g7
E1:_SH9T.YH:KO>YTZb9U<KC4_79T5P[K#7QVP&S7H1KWXQ(<0@:HF.f5-9/JEO\
<K8H)U[+?FgbN:cV0&YX/AITJ5WH1OTM:+AQ5/gDM&5[DZW:c2aK)AI9GR)BKYUF
/-W^+=aeGX57#DE1I+\\K&_a[98.FNK\IQ^<UD)VR(B&?#F@M4eGWO&B2ZZ>Q]&L
S.7PY6Fc<_NGgR(K#0a\GZgYT0?K9/\=)69VZ>JgK0/V#C6K=;a=TZ:(:A+4/2P^
ID6<.61<TPG8KXgdXS3:P.<1UR4>?eN>[&KE:dOdKHYT?GZLVXZ?_]1E#d#V.>&K
?a^gRW++900;F22H&GT.9P:5[&eZ.&JFL\D[224(fE\@WHN[46=XcEET/4M=O9U>
/g-I=>QHNWO;aO\.f0RGU2?]@GK+&[418T/S38K#JVZ\M(R,B4DZRQegP=99HXc>
Y=,g()N1Z>_@]7.XA#WP+Cb)^Y)89gU^CHfbJI:&AFJ9RH,D?BAbI2RIR-^BcU&?
[:afV1RDX1JD0@-HF/F#D7RYBN\S32L\Z<M#?7]2d-bR_&.AR6.SU\,50\dg-a6H
8TRLcC83C5.ET8089e659+Mf</\6@gef]4TbXYb8cT3+&#N[O:V5B?;L;RYW+O^/
3CaLTgGXfZUG6&D<T#DOHYeW^9;G8(ce[SR:5/7B+9&X>cP(Pc5e?aL<\bAPJCe1
&5g?b(B[[bN/^69LOI6H6?RQ51P36,IT@F2UHBSCPf]I<;DNX8Q+?5?Y1Ne;9RW<
-K8.VS5QJMRJMYZ)W9=Ue]T[Z1VV?2(O&VPb8X=c<-:#&0g9[>T<KG0aD)L_?fHf
IS3S9_<_[:1aD<U.YCUNY0=<dfG52.=R2WHE\d5MFFB-7D_Uc?1N-(Y:MMI(IOX)
29?(5J]fa\LC8#>F.6GIG>OePD#32fR^MTZbVJ.(=G_.V6>7KWCQFaU3@>3Q\E(]
6+ZNCW-D0aA6c?fUOX96<b#2gg6FE&8GgAS1.bd.-A:[/1+5PO=5]X79&G<\Y[2&
U,UfJAcC/3d5Ae@V<>T.TY6fP5R)06F/BED)NW8<<BTWIe3<Q:.fSR:80P.@DODY
U#+=63SN8Z#H2c.81+&(X;D7;VTcQ2ae9V#Ua#QUKJ-98cT#QA&&LA?e9:P9bO?:
O,]9?C@@_=KWYTDeI9]Oc?)(S_[69<HU(=G:LQN-I>?E<+bHT0,[A>RH)JOMDD?+
U_QZB:WdK)[AY#)&[fH?H\e(J[)2QTZ:<R:QX&E7JL@]-Ha^XPb1.)/J_#Hed<)8
J3f6J9)AHc2>21;U.16#Pd4R<A6Xg:80]feYFV#8:@Y.]#G1DU,U2.S8dOg9<&B(
fHeK@@G/<c56D>5LG+9N7;2&O8QX/6D@]:JWId\2>B:./&SA]Qg9BSYZ4M(<8&-a
>Y;-/-\X1X7B_ET3VFZAQ<&Y&4(I_6W[#VCUYb4UAef)e\f+24G:QR8cS>_=X#f[
FBa6#V:dBaScW;)&._c119A#88ZQc+?S+CZK+&Fd>WNQ)b1NR1/GGX6]#0F=ZZ9U
3Qfb)/]7(]MRICSV@WAc3RD@IE:L\g9UIDXdK.Ngbcf@HD(PRWORL\?b[FT_H;14
LebA8&ZPK#=QSC?QW2RMRg:UGF_^#Y89^\VaA]/;fda]H4.Qb/g,4-(_;(_KY@eV
<4fC8](>JTg=31CF+&SYEFRHC5RB#E]E&B->CN>IC=3B>I>4[_2,3g.=N^bZO9C_
//#B#gL#&L>:_E<NaO\\4PYI[4;2;KE=Mg8GO1DR,W--[R&^HMIG,D429QBJGY@T
b^a02).2_#WXX2EVSRD0H,Fd8.c&FO+DJ/G\1>P9,gIfN)KW1LdJUbE#U-#=:a6W
BU1HWC8&=]CCc:1)Y#Y\gbPdA@0NVA_\J4<^X[>D+XLddHUA6eY[&5O3TS/.-AU6
]SRTG77C(dI>_KTgQXAbR[2S5AK147T&&XT=DI.LEK,gWggERPV&LSIRS\9GBVFQ
J+0_AF\GO&^9J]C/VDZ(37-3&KVYa=V&FMJ-^?CIJR.G/IW8]1]1>b5QbPd.HT.=
8VdOEH@fb-OT7L[I;X0GT8A>S#PJ1dFWC)SZHY_5F.YLeL4Sa<&N3F\<#^C2&fV]
](SF:=X&#F7]&1SRC1D;8b:8&&0=BCMI)6>CS4YLU@H&dNbRcR_QEVg1YG4b=L&U
#Sf#WMgGSD[7dGWO#NL;J&X4c)W[67&VUU?&:?2(L2C@:Ha-CP@6cQD_/V->;(,@
[RU-U3QSQg:U.e<P927,D6ZQ.bO7\H-)W=^:+/fP/&6fME]ZBbJN_G>\L;YL/<0P
f&8V@;2:B&C&-c>:E\T;:S=Be^[:7/JKZSdb;\Y.XUX3SIX3O5P;0.DfZR)/c[.^
XKGN^S8E)0;C@GK>906,U#9LIaB;64W5eC^U03I]T=MdaGK5R<N4_&[E<W)9S-QL
PIfT473P>g@/.c<8OJBC7_4@]Q>.BbEd^,&(^SJ^@7>@Yf2T77S9S<?__5TXcB.I
2C>:fP@@7#dGHcCfA@\?:I6/=>]HVHMKCEaH5D.-ba^;TC:S#UOC;A<\=/277X#I
PfSY?C+.H@BTT6I9A8R;V3]gT;c@4?LYSE7N,G=&c,19^UNae7E0#]/(,6D;?52G
U@2^EgM^P(QHdfS(/ge,UMUKVM1@/=.67eJeDHccfa6ILE92N6]JeGF7#_.[A41I
42&7N#@E66GRFYUYEXV-<X@M(Q.MW]K1Fg\U^Vc<:3-._Q4,H:8POMBCRLA5OI3=
\OBXRSAV^T0a6(3LB&EY?1KURD[]3&1)14EAYDMM>Z#IQP_8I5eMT\=V+]Y_fL_\
^WgN/91?\^),&682JWF\(>gaFS9<&.>8_6+5?TRcI1bG_gWRLTTYA[::@eL_+aeT
7+R(cg]A:^+A,d7RG\9;G>ILbABa6g-a<#^E[(\)>(OCT=Y#VESW4883#7YSX6VX
P9G6.TX2@L;cID)YHK[,?#e_EA7]U(5PCNO&Q2IJ8@KBV_C<,0_(DMC896<7<(:5
L>Z^6OYWN3&Hc3T-+0SGUZg=,aOA+W\/H=<84@U<B6_7g-JVN1O0\O8O[<966.Y,
gbU/=6XG/?RAe^)9cLI+:75.7P4M;JRUY3gC4Q\KXdc/dD..#1E8_84#J;-b;K--
UF&&cBPgVH4BB>K[)VE#J,C6_cM8=P:3Ne>H>1&+aMaGS=XfLB#,AG@9dc,;Na4X
Be[TG.8[SP(JVZ]/_AQ>YPRA&gIY=-<J-d=ebA[0b8)733=RH<&.&6+b&0<[E\S+
T=@-)(1B096Hb+MM6O<dDKL]IQKJGeQT7ES>.FBGU.^>R^.[c]F/;E&KL?(aJ/-U
MTYc5(42W-[1@&RE,Z@P11O])56I&?,8\QKC.9IcZ)RDMLZGfXJT0YQaG1IGCJOX
ZK_PN\C:9,fFO48Y09&#W>)?-.WZ/9gUfUb+gF]?#D?N^FR.]JRUcf]GADg^dcVg
NM84#_H.F6^EPME9/2OUgH3:W\-^A-D.P@gJDYT.aOAaS27X_/gCPVCVeW]OUK2\
RT\6]7d3,7MWBg_J47J^g2?U7\8D7D6SNJ#)[#+:]\D.b&]:1A0?CC6)Gf=IFOe.
K^Q7WB.AQM46_XPeW.Z;a747>b0S6QJB<6RPgKO;?eT#[]fMR]:F>aV)@]]UOJ0<
N_;BfPa_UW;)9S..Ta/c@-X4?aA?+1B+4W3Fa3KMU>><BA<[8_FZee5.<L^>3Z5^
=+I(3AD#\SAHFbSMbLX+?B7W<FJ@)<5QQ10P2FA;LS(FA]W#/2RM5#].6E?W1[)A
7]\NU=eKb)O#BN4gg#Z:0]YXAWeca=?@<LCT4<aQb]IL,c(<H-@Wb]H^LL9Q@)X-
_&+[f)@eE/g;TIEc&E8KV2NB&dUd/+GOSbW):B2]AGO_+#d^7262K2KM1e#:e^H?
<=H4@[2XH&::L(X.6YB1SS6MZQ^[BSf?4e57E#e3?>Lfcc3IZdPFaI4GA>]W<cL>
G(B^+=BS?Ud;2fL+&FP&YT(DQ+Q>dE@fE8._@H22H>UZ0:R9,2ZaLe:U[cHPAQ[2
3,&\f0-]TL@66#UV<HP#XMT/]X+]-CGS,.MfB>ZeEFL/Y)&.V17NT-6VRXW),c#W
-A&FBLLARYXWDb\Vc07E>FFQcL,2#0>V5AO_@N8^VZY(2:HJEI#RB\LPA7QK<b)J
/7XLC#8+[#VgUZ[Y5Q071P38Nd4cKCV=@Y#95U/fe\Z)GN@7^S6#7/I-B1=5\WeF
Kf<VFQ+aebA.<-.;BR<7?gc/b]9Z^HGG:.=MYc^.ON72a_L[3H1_3b[aC^]-(ZVZ
/;<+T#_6,S>]C.#5d675+/O+FH9GBH-7+?g0g@?ISQ;MaaTb1B:/>YZ4=V5T@+4.
bQ]N#HV=Pa1,3?K_N?cD_4V6SKR[6(cD\Se>fT3Gd1UGM[cVPDb+fL)KD?[^[-5^
E5dKSd;>OWg>;?S<V/2YCF9?F2>>=4,@A;O.HZG0?OD=K?X>A2/DW;1372@_E5PD
gI[)dZ,AI)eF_NX>0LZWULJHDF1I5FS1^C6<(g#;]+&fCKE\M5:6g7D[<8&),7J7
HaK#gb81d(_[4._\+5VQ70D3ZQG8SEE[TT-5P(2Xa+OO],a2MJcBDZ,_N@8K>-MM
QW>A<JX(Y0]^aCPYDX&77@_ROLV=/:>C_\WL3+e>VB7^8_1_)N>a<T0<WBE@L?<P
KMZdJLc?WbJDU1gf,(U<f\IE.-aLJ>1f5b<XU,V=IELggY4f:-[dLZL\)L?NP[]P
V[43/1Z0>DPG&[CO.R=3bXTQT0\P(D8aB\9#QBD9EU=>AED02F[H\ME<TP5(SO8E
1&\NQX4J&C>5-UUN_OY;^?H7U>GE0XMM5XS7Jf0D=(#+X><1<b&(\V94]VPd:5MK
f/O=A9A2XB^&E&#>5GHPD;QO&D+,g;Q(D4VR(]\-KWC^6ZOND<YQN\4Ab8EaQd27
=<ca(P)B-?6b095N.RJJ)NFC0),^F))1BV&b.21H2[/&(F+RL;YcV+Ng#AK;d1gS
8FJYNY\3fTM8aP1,A7<)GDX:.A2>1^R)1eK_,Z)4PC-KKJ++R5,:19SbC>9NS_NW
+,>e@0RVS:.;S?TGWD>1<RQS5eN2QfN-7_Y+MM5\7.3SaFc5-J<\#0<@J2?-^Gf&
G^-<KTN;M[Je6B_([KC=\][H1Ma\-d#:Pf?S3G=V^<?2Q]^?-[3bc)?.NXQNfB[V
RT]EIH-^J8JN-ECRS(7#I4;][?S(^Y-bB4I8UA]dVBa&fL_f\gW(Hd;UT);&\a)Z
B9]D0PWQ#CV??4AIK&0#M_LH,G=_V-8.?_XXeI62(Ra2-D&[BCB/V=X(\06C77g&
MQ68SL?M:ISF^E#ONQ-TMB=cA_R.CV+Z?T5J3NC6KSNLa5&c#(62I>=PEbf2#FQK
W?/G^@[Xd8-MTHT(1VC8A,a1++&=K--),HV,6D<eQCKN0&3UFSK0JbGQ\0FX-FSe
7,-e)XZQCE8[g;fVA/H&/OEU;;9@E:D0M6#-9_f3V,Ua&9.8M1>g5+J,QNT_3EE0
G7D#I>0_#Rga&g0;ZK==5I9VENA+P+^/-2NV?2AP6G7Z+GR;CcHc33.KA\AS=QES
8H8\C9c@N)IK1M>V4c76G^6@O2NA>5&4[\V4PUAf,GXPNJaCPd+S:Y-MUV:M#C4O
BNBP<G[N#IGRcN;dV.W+A:T,DaZ.9cOG^/)P]@O>_b<KA,bHa?4S-QY3e/7T&DE+
CG0GMe93N@=@.DWVfU+--C2W@.MbP=<Q])H<;G)U[dR0MJ9IWH0#_TIV15LC:aE(
U2?;+5^7\28Ea[2ec^27-eSR3aYJY)4-#WH)FJY)9Y,4,D/>:I0@8KGA8V1=D+[#
Z6f_35LM1I,dQUf^W;.6<f5&EG3@Q?:-)U&#UB1#?&[O:d2O2YU^OU4Kd1Q5c_9c
<#d;#1a69=@?Z8D?AON1]_3c)#,Ya9R<@2?gXff2RSc1)e[DT<50TgJa?fMY@CbZ
7,@67g\ML\R\OS1B:g2db;/.D@<-,J6-F,#)C?>.c=(=0=/G\&5(&TgNdYgK;\8=
07F6UGgH9G[JQKN&5C;>0WZ214M1E8cRA/Ife8]#[2J=G]:3&QWY6DNbDc&A?<JB
A+Z/cH#b1_UJHV==.1ReM7T3QW:.7)7(DT99SD56Gb-N8g?#&,:N#QS>?e3Z;?Xd
:8\V9J.b5MP=>YQ4<8XW?Y]4O&@DCcF,7b?.@N0+d-1Y^LeV,3H]WL_,a1>/.QNL
[B1aH8#[7-MP0F;98Bf/@#N=3N0O^QBN@S5dEN^3IE+<C8.1FU?0+1I:NZUA[7Z/
3g,e<T[:4:VZK&3gT.O&UQBT(CgPPDT-SFHE0O?GBI[L<KR@@[?76f6]D7?+?+6Z
Cg4aAEW:cZPaTF?(+4ZI2]dT>GW)89F[SS.<WBbCSL2+M.31b6Y3-]@J_;/dd\aI
#c-O?CE).J](-6:CM_ceAdLF9Ldg)T#E(CO/?eXD8W?WWXEZ#&7+Kc.7F>b^2\L>
IXQ8QgKH.N8QQe)L[GJT4JPe:IXB<cNVMHdLFfTga9\^GIQ1G^d,c<LT0bdP=F+C
H=YN:J/8f_#.6W#PLCF0X[J6=Ke/bgM,6HaM9IXbZEc&#W<WY_H\>D3)(\/]3:=,
PdEQ#EP2fI-,:c2,DFK],9<SUS>UP^)G6KA9\fbX\H@7NMQWPd=LcEAEfR3R\/(Z
H=UaHb_,PKIRK4I_NH44R?5:_N#0&#IBCI?G,9Kbc[@[LdL=8VRJ)bEd0#:\K5B1
0K5T:E<+NIK.9EAM6XHX]E4aBF);]9JP0,DC+RZ>c\Y\R,GE<RDc?OM1>,/(4K>]
Yf,I>5(c-bOR(aYWJf;PL.PTKD[GLMAR;W,#<XR.HgJXR\RU7?c;ODA9/1Q8>.a8
DPOOf:=5eR6>+68],dc3UbP_GO1\XPC:3TTH>SI[<8C8.D8)b^8Z(a5d:Dg:1S)@
+fUTb/(BQ(b5+GIHW?UUU,B5P^?->PB;#J(D/UZ/_I1F>^/.a;K0,Ga/KO5P1T5<
9g[U4#./\Q<SQ^4L&33f38Y6KOA^.;3=9]Q8/9-0e0TZP\2IJ8:cV9YJY32a(P(&
SbWXb:7.KM]Z-S&;UPTR.800#FZYOP@&]R&C/@]6B0K9+<5[<4GP,,?g=5S2GW1@
U_OM;dKV=N1db4@(]g#DQYZ,R:J/T0E\Id[3]cFU4J>7KB0AIK2fOBcHI3-PGV7M
S1_LKNd/+<F5;YV)B/;Z1P-JaWSR&WQb+a_(BeDJ.MV4Td0V2X3OV5:a#.Pa@_A_
,3^&\OJR:TFBFc_8Vc^7Q&T/eD([XMNTAIX4e=-g3:=eX-W/#-ScK^_+W@B6C2A&
PVK[:5Mf3a]=9XU@-U4FF+1)P23SB>fZ6_]^OCc]3>^<FDdW81@^DD[\;W9([MY7
3d^RA2H77EQTI]b[bf38+]#I&\fg26G:[2GXM0^8-,21&8CI/RM\>c>N(+:W[VBA
C0.6/cgC^77BKQ=2=.YN0]8YK3@:^N:If39E&T&E0f/G^+?fX=-;]Ra[0SQ_VP9Q
2+0V_5(g0^@D1\=P1W^?/G>+3L&V4FHV8>fN:XW2L]BV2RJMLF32,e_g.X9TZa4)
Ma;2MFC3=J<BW.b_1^_fQB69@Q0AT/(TD0&S1&7,@MAe?e-O=bE-Jgc8-S35C4QQ
B]^B-.K0HaS05L,X0+deZd^=1@L0_8Jd<BNE-6Y_V<7e;_.^Y2:6dNA.&W)JaP^/
-2KEVaZXZ?MLX\JY867DHdWV2c:AN2=(=XTLdMfNE+I7aJ0fLd9OEZc/b5,O470C
A^cf]YE;dcL#H7:K59:#<X2<0#&3;[97\^0/_2XSMKeJ7PKd<9TEVLX5.>BV?FXR
^CB2aV_Bg1S-@UZcf+V(MX#W1S_5XgfTE?-dH\.g/dWSP7:M;U\ZCD\E8Z67EMd=
#[M6E(b@:G:&8f2#^[a9LfWZ\[3OaZ6H^JK5]9]0LE)KGdFEKG.Ad=V4_5KLa9:b
P>6]-I,(N,9>BUEXMN>U5c>[9cUAc@Sg+?N<=2D_G1_c>>]9SZgE@50_=M,g]J.H
baV2@_ESP0(7#:6P>]DJ2+7-bf#R763T)8KIZP.W.#MALfB,HOAE<?M>A^#KIBDZ
A>7_gbK,Ib..9G9NXfCWJ/1SVf6&41+OT@FR&>^CRCT<V_LO3Md5_QLQTX_1C0Z_
5IaIZQa](0Q;g/^GI-ST80:?e(AB,0f-R)\VAMDb&gb9KD?@D]c?FX5W555F[a0g
Y:Z.eF82GWICfC@e[+BDKIYT.HPg4,?[J[80W7SG-J2(-\ab4#04&]CM8[J,g[(P
Q<&RA:;f0cVMdR5_dPLT_9BYB^1bZ4DegOgAI^^(fdV0MNYJ>[C;&UJ;(6FS17cY
UT>_=C,L/9-_&)(=6D=AQa:W=5.G[@WOZC2@=RWOYD=#I8a#0eDY0BNO6bH<Y48Q
[+_V/#_V:+#ZN2+59G+WRePe(eT^fO-?FVD8D0TEJdS+1X91H[N6/TdeW]?Y,Ya5
;bO4@?R=6EUHB(K^cd1<a&NN\SK8II>YE_4g<>bKC=OL&=,@c)H=Lg=L)HJ.L^[9
3II2K7/_Z^.L9I6e8/J@]f<A(>5HSM[CD/)N1+>Z5VZ7g.1-bV-GOK+D,9=#:)W_
WF>IY+eQI;g1gXJ1Y9f8E?<\U<eQXO2P:Q=(UK\&J0TKQUKNb):PQ[BZ>A19B#\@
9CQ,8E#D.FI--XN/CEg2RPAI>/)d04Vc2Y@J[-W\)R3E53b<f-3(HIONXF._.acY
HEc#eb)OFLP6B&V/+NDH>D[#L(;>.&.C=d);a?4Z?W>KA1c^EY#E-+2KEI];=>5R
.g_WcM>()F@I-bC5]cU0AH/@A;P\SBS7fgK]_,D>\VHO:(gdaV7J\Y)B=?1\B+If
XDR2+gH[;Cf(8W:R]40_&RSBEeA-.VgYc0TK8NOL[-OQ;&Z-U)bQR?>[>C(^O9Of
&b0ZP74F]J/4S7]WG1Ed?fYaQ[)FDLCQ5@A48H#-7+>R6Ef^g&EP^@b9b-(1&3II
NS_D]LCKS-fe[(J/d>_bRG/L[4><OG8ZD9g_A#D<E0-W-.=.B40(S=5KIaQbeH?d
MV\GI<]_gg5_N76KK,-D&08W2]Ng=;8d\#gaeWJ;=PMP]]S5FVZe7gg<6(N+):(R
PV&X08Yf4W0]M30^/@=RL:Oe:BTPO&fe<,#bRME<d;&N3Z#AK6f7ag6C(d&EK8M&
WL3T7+Q8G.,3<ZNQQ]SeI(:W^B+W<RO2dc>g4\+H4Le&T+N^>27LUEW=5LgZbQVF
IRL4UJ3T_W0,9.3L,+#AY&E,&FUaeW?B8.KPG9&Lab;J[BUd2>b:Y[5W(/2E--DT
04D_7_a10V?Y)M?Z.Yg:D.]H=C;LaA8QBEW\)4X]\L@M(YFH3GF9RP@/L;Z4RT9B
BJbA7\S6OQBLQWP(J(M2dG6_PR9(I2fO.>#GE]c5GYYIc41:Vg/+[.?,8/>gc^W<
g(Y4I0@@T4+1CUNH)C6T?N@9,=B\<Z#a-C\?9Y==JUI-=QbfYd:ec9L<?H>3.XI<
Q6#J>7F?4.<e>P\>HFD050:2N?G(WSINA<R(;DH&cM,aY-MHg24(DA8D7<A5#-K?
c&YX4fIDbVRfB/:ZIF6T@CHg7AgY)>G?(e;df&D[99+#NSBW-\F(e-TfLQL(aD@0
-].;6)^X+<=DM.33/M[O10E>X806=Mg;Zf[(Ta4IKA6H#S^@/Ig_NS/6d\;.<@3.
P>c3FXE()BV0KTN3HB+?YCTT:cca[FN-EE\UT(fWZYYA\H_Sb4_DMb&,d-(G@\^G
X5B\VPQHfMBT@\L\^dRS<SSY[SYT/A\)UQbLF5LS,F(7e]#>_3\&=22C@Jg(GgZc
+_:9.G8DWb67PaG08+5+Uae1G,YUEHa[)@M@]S,]E6(gL9]+Q+U7L8MLaY2UZYH1
R00WaD(-P8))QaTL^#PN/bIO36aZ5UKF&&-9N?#Q><X2W=c<b;)(KcbJ^N-Ogg^F
YI858C)WaWW>fK?T[ZE^)@]Q51QMT,RBAZD]0X[Q,ZXb3b]249[(5V\9CeT0PHRH
eBYcKK3gFQWI4c)5F73ZX&+Fb/OXNEC]0]?[I@1?&#cPE&gN-1TK#7(PbS?FT:S=
9e>8O[Ga8L2=ID\7XCg_XVU#G#][Q1G3g^>A;CKTeZ@B5+QMM]<0;TZB0KV^-XV1
B>,AF?TM;FeL&M,eDNPI>P&ZB59[QdGI-4PS,9A@Cg]Hdd:65=+c<SF]M/L&,+12
D,9_+2,bUf8)\#J3&8Hd/\57MIZQ^S?.,>fGc^K7XD)8K?g?/ZXWAe7LNMfbXdT\
d35<U1LRNX&IWg,X#9Y_9&#WfQK>;Uc3NW>XT[,L7(AfB,LQAZ<[0,D8cJ-HTfE0
KR.I1W_GHAJ=\MQcB5^=W28N0MY2c&8:cM:^))OEHR?#<[Z2=M?aU<bgId-L@5/?
M-&X3@bc;U-<1RM/<,<R9._=aHBgAP>4IH?7A?a\?1d<g]]e>QQGaUDc.4fY#[))
OH9Af)BE\73&;@]:5^P4,[X<T\K:BVZ?ccTbCRU;>>[1&0P-:5b0UJ]f]6bff7VV
P9&/_?E/)NRG:Zf[6G1&O6-+&(#21,YcF_+BV6[fS>]+KD[:])9DN#A-1#>T^P-;
7UgWG.]C)>bfFWVE+0dZD2D;eO@469@K@DVZGf)(26@V>+6]>]XO8=N-B_GA&b70
];/F01HJ)KUF4G3RIKI\]K,]GHQV[#W:MT\2:835;Q;<J=R0D2W=M7GB)Tec_+F5
=S=IUPgJ?FfN1E1F:SO(/,ebD#Y(2)5J5aHZS#^P9X9RBNT)#f(eL?#XWHa^fg:5
eV#NXZGTYD6-I,XB-1b)d[79,;HWO3/?dCA8(\fJ9,UWa)QJ_D(4<94_N2]a?F.:
?N<5#Y[daRZeR<C4YW.GS&M,cbL9P#Z<FXf3>)aTfK2MfcG^NFZ/+8UK&:V,]P?[
]/O4U]=7Kf_BbGKNa>./Y?N/O?c65d^g(TT@Z:eM4++:W:M@+1+>&+Q3E+eNL<#D
c3<47M,+f9g1],R_e_TS);[a3-_HGF1M3X;J-b_P30],?TU_62OSd??dRE(8CV3>
HWE2c)O#UQAVUf566Gd2FOQ2AfC:6<eNH3aeN20f:g7UgHGH,EC;7OB?H3@&7F6M
Z^S9]?Gb)7L8NH202OA?c1#IX,D/eZP+N))1NQ1BKIII/NO:PabWOYb),)0dR3-0
A-2f1;:?W0CQ+Ub6]L#HTYRYI2SF[]@edK[7-G2[RHQ/5Z0MfVdBI3dQH[1MXa[9
f(/NUN8[WSLbeXJDAU=D2dTf]?.6OL(00TR>0?_N9<@:Vc8&]KZAV?gX&UV[ATD#
g88f3eb:GE;ZAa6D>UHHNdg[De-(7+#W;bO[R<3Ede)D0cR9JG@BHX[E[eK4Q>PE
@Xd)@g-JHL^1W[f]>@#[<ST8#,U<?95419c5@+a?@eH/#2KKM1BJWH[NP3aH@^<C
&+]ZJRd6B:VAgYZcGZNdPf3F]F(P#?WGPYL4M7R2PP60DA^aFKM?+O#YCgVI7_[.
7U3gS.0DEJZ.),^bCDLNV3#GZ1-(gQG5J:\(]X=#,U,CD?WS,dQacbW41a)QI8a:
ggSLX\7LA.ZZ0c;=G2UCJA+eDHeEJHZULUIZH0S/2B78^KR-e)6Ie5EL]_S6HMGP
S0MB+c/U@D^+8TcD5ZY9CP[X(/7Z8XULdPW.5U_@G_@OeA1B?P\N,FZ2A[dP#[V.
R-&9JKH;_OM>FBgdJ_LBX]=QH?P<FK8L2P1]&gN37^VUC.g#(Gg/2U(UNTGg6T:a
HcZA+T@g#.+C8B@[</D^?[fba3VC)F8)AHWAGU+GN3U-cY\JAV9C8\IZUb=\Z^,R
7]82]:P1;,Aga\V7&V=XeUebJ7IULA/QfG7>_)T;>M]+Ec/7+=Zg87<a0#>OZg,8
Z3eY3\O?)(2;ZU^^RO,8@;AX\DCP6LD?,-]b+B,efa^2[>),1Jf;VGBEQ@US&O5C
C1dM@M@R+Rf2K#NQ\HW8<(7I+WB[W48TfD4fIKWC[WJ@RF\XGI<?CbDJaBb4SGf#
\+b-UYZDe2@]_NYffU_aY=A<B3[a>=98GFHVNfTM?Q-3(cC[AJW:<JOd5a0RS&D;
2Zb;D:)4R[b;\JB0LaHH#=N4TRU8S2:;B/Q(Q_#3<,G]J[QK7=QU^TE]b,]8;3O@
7EeJZTgXXM=S#:J.1P@>C:M3CY1<,W#MMQAQ93)G\^^=[8[LUXN1dIH3U]Z,/2/A
:.C#cONU(dS?&M-<35?&H<]X:,YT:NQ1,&5YZ^\PBO-7&::cV4E>)MMUJdeW9F<]
GJbbJK=VN1DR]+UEQW[@>N(L&3#HRdWZ1A^_DK#ag8U<0Q_-a>d+UMV^[+)_4/BX
24YIJ17BeD-KMDP+g(<C99)RSA\<AJB0c5>K_\/KeM@DGH)PR[[MTJ]X^[&,NIgV
beWX2]S[CPA93aI^\25_2,:88ZR8fb^4&>RLdbX0V#[\B9-JV(\SaR-9F<Id2I8W
\ZXJ,OOZGDRT=9[013\dQ\[geJ;+#[.FRK<)_G41RTC7-(Kb)Dd;Z(BgFYX8C&53
c/.g#DW5RU\>AVXX=U4?^+UO:UK&TPZ>R\#6@+V7M1gG5BdEY??c-7??2T=:bUaN
5NKS&D]>7<.a>4dEW/2F3>PeX@THD;cPL@aV=^DFUP^#NO4Z.SKFQcd6OC@#JKbe
Y;A\_,0)Y>28TC(->]:[WBcQGgA?b.MT.;=\FKd8Ee]d_#4c5R,<I.f2+HDaALHM
H3-U6USOL)B2\d1^#C.#KFNS+_a52H.,XBf?T7^Ig=9H9bQ2SDbMM8_99)0fC\CB
PFLK8fY3/PO;^&<c4TGOM]S^Q0GKTefYdQe9]LU>gQIH3McP:S8(BF4.V//#QdcN
;[=<a(I/S1:OW0]8Jd=Y-&W;Mc90\9Be?/#,76F<WQGaT??C4_J1R@fdD_/[0Q/8
:eV?X7CH[g27>HV?BfDAAN6a[UN^1#fDL<;8RGR?LSQa&>b6[0CMRQ_DXXfZU5aA
DPMR:dGW.0(RaU>.Td>2)bc6NQ,f&THe.NW0#Z#C,fb/I5TZPK(W,YZf8aPHZZCb
#\+Z84N^BII9Lb;LG1YQ1MLD9UM<?VO3<L-\2]a7PGb6B-_)U:FVeQ/>[50P4=PJ
;QVI1LI4g.g8Nc>]bT&ZE>##B;AU1;0IT\L1LGB&a1M[J24>1537)fTfZA4RZV2_
=d]ITD&=:g&\DSHUbff\O4C;69)6(89QSHJKGCd.1:59VO]D_e?7ZGR&R]>feTBL
?Xa(a^TJUMUXX,5HD)3M8A(C;,1XV/IRG/2/V@DOe6H)^[DL.M>eGWH[1T6?7@83
JcN5?<F+&Bc;>(CgIS#\0>:?)H7M<^,VOM&g^\T@,aJM:CZYf5F+BZ9>>M61X2N4
M73^S8g+Z\\OY;7>c8?HGEVd#];RGIQ37dYY>5JQQO+gaX6&^17JT?TW5YeVJQ]4
C;1EgHFF@F]BV#+F4a;U-F+R>3;U-1/gN5K?>,]A+Hb@GbN+:3-PNK5MJ;Q+R^WD
NU9V=X\F778CX>E>20#aLgFXg<Qa\#O[554S(^+beC>=77a_S);;OXT+VTIe6@eN
MT<#XeZ4ZFeedc^bSW4[#g+Gc9[HB<61SO.[Sa?]OdU)G2Y\9#-e-?YMd]5caaIP
DO/Ha)E<Tg2Q,dY]D:P<R0R6UP<bY,0;:OS[)I[];K4/13L4YGGTUPDWE>F:c,=1
=QFG8Te/d.+A+[;^c0cXB_D(X#AU\cTa5V>\WY9gOB_AKPL..K<gS;g-4-+V4<AD
QD,3##8@]&]DRgR?L-SPGNbEB1=T0dP^=bI,)?Z]209G<^2T=b53Sa:/;,_F6@dY
?:HGENgf/[X5&Z)R&8?<[;(f<.UT)(+^(M(9()L?9A;.D,AJdVM./9IWBBIU:X9X
g3GV+EMX2F14?7R:(,1-O)2>T^(=DN^eKAY_<#DfC5\VZ[G=_VOeKCAU[;d)Y.SI
c;,0?ZYg?0DeaRY,WW)-QS:DQ4>LLCd+\^8a0OZKH^L+124#\.8A+B/L>RMYIS&M
2_Zd#Lf<:XAMW7dS14f=g+3GK8ZL/f(WP_;V&R@eAUF_P_.KN\<#\+):,NONOaec
M>W2_[SDNEHG,gZHCeJ/AMPFU&@9+POKB1;XIJC]VV:N[eRI<PQb/-V:?\B&3NA.
)EXWU.0)T>&263eH4VH2&8@>(]LF?^JOBY<VWW3[.?HE29eJUG<aGc4M^[/XT046
6+3(S#]Q.R^&VC^B[<?(Yd[gL.)(),5N8,LK+<KNAfMT&EeMQQ/\#BH0F2D+.ZCN
Fb?R4<O4CXCc(>=0f_I52bI[aVN?Q@D(UD0&BF-61db8B)DZ6E<aS,@fSWX5[J2)
IPgFYD8MIUAg3[1,>B9[8g/K?(PS:41g=:(T^+0[WG_BN^&VeaL->D)64HAI0BgQ
:a-@c:XgcCR&@EBMPIS82N6WE]Y,dfe<J_5IE&.aZP@VGD-a_c(;JS2IY?J9[5IF
D40O(LEH]R,#SZWDX9,&AggOOY3F>>0Z7](\EUOcd3=+^L+_&(NZWHOPZWKF4ZXI
SW0>:/R3K)))7FaX5OLS8WI1E?3?K.XNIg<&6QUTM<&V&U(CS[HI^9VeA=eVcQ#9
[03D1C]J1V:@&HL8-e85_Qf&8A1QTA3c>Y/YQcS#ZH=IM89;C.9B:]CQTa?ZDE0#
YFM+GM&R+g=Re5Ad<=STFU:d(D]]D0S)H<4&A,#.Nf^DQ(3[]YgKK6f:JX-0P0FP
()0\Z1MH5OF#e7[dJW92-\Z^8A^(>MS=>=/R;KXG-eg6K,d5YZN&<5NJ[09EF0:G
<U1MbENBLI4gT9#M\(Z;P/B;]V,GS,C-7X2Ob+KJdaD4^J7YV@7=9BATC#;-2-GU
JY@OBTLfAG,>/Xc0(K(J\-7?^(S8fDP_M+P&]cK;c?/N_>dB)Ec.4<1C4Y.&WT2X
NVUb<b5Q,]VMDb2#[/=eU<JHa[&6;]4YMg<.)][WR:UAfVIR@84D0]MMRNF1J3a_
E>bO;#77=>-5>H\576+eX(DOQ-079O4@MbMT14M<OEPOCE7UVc><RN_E35L.2g5#
B6ESWW_B#DB>S/7K9c<e?[U1\9,KL\4J](+^ZS#MUeOO_/[Q1K>GQ-7#YN@>2V3X
(O_eeXKF9a_L[EXSP8gL&c5AX)>E_/NP5JAJ];Q;cfg@/bBKFA2L<g9a1+[84KX.
+6&Zd?NC#NeS\Z-H3fOPQYcIe.Y&P@GI1BCS3+&/ZQ6Z[,Xg0eeS(\Z51bOd^PJd
:(Z]&MM\R7&6Y8Z&W=4,E:3Y&0B?Od6/M.Q?K&05;,@CQ/]gJ:C3KTfbc9T5QQ9(
0Ld:D16MHQHLd-)fC.@8:)?V2J<XARO^KLKL7,U9b>?I>[SVVE+bF.#WBN4#9D3_
21BW^+9-8:\f?SU>9EN?COG9[>cgc?9HgI0W;HRgB(->aSR/[,TB:[<ISf)+#ed+
\a:_B0]?^</cR:>B?^F>eN;/1;M0<UCO?Xd\J+?6P&Be+6QO:M7C[(#f^K]-S5C:
]&ZT80PNG/7b6GU+-,c9D<KBHBF3(<1-D\G)(5U?4GC7H@P=JWZ7=UgJ>aM;(@KC
]2B3>^3(A^62Z?5T1A;VPN2V94bK\0]1YS33:A,c@>YE+5QRQM;\-C@U#G?<JS?E
?-ddEGQJ74.1)?]HCST;FAGX7:KI5N6KLPa[\NdO(g:[7H-^&\RF[e2>:HNE]BF]
\L1ISOIdaBPC@bLX.8=32#9A2R6K:4G=T?4HFc>X5Gc?DQMU9dIR@>MHW1_7^WB+
XC:@@)Q1e1@,bN][N^MY21c(SUY/O6bXa9N?@IWdZF3gZfU;c2?#daJ?LbcRda0_
U364JQ_eTG94A7-aYRSY11YdE-59DM<Q8Y9/]2?.P^HJKT/DT23c+N/ARCaTRP-C
(;Y,d.^]QS7WB=;:);F@D6&A7Qc]B=^OYI]KJITaA0AT-Z?>V^I]Bc68<^d9RH@9
\;/9LD/2]W74Tg5H#/\0B;=X+a2.?FdA]0,X(J/G3(^FGNK,H,PIX8.@W903Y69g
]@>7bcH-2QE94eT<L+8>R/&21E1eQY(K<H-+8UO7R4f>eA\.CM(U:<(f3Y0(;d=W
Vg[UIU&?[81e=5X[S638/U)ZBScI8O#cMaPI+0;D?XY?L?4QFU>[+fMT+1YPI3_=
3BS0(C[II,<H(6@FcM_aYTQI[?#H3PZ.YW&PB^SSb:ALW7[G1\S72NJ(15^K[8#N
/EPT_eN2,+Ag<^fXdKKT,8R:9QYDPH42/QJ4>@:<N07Z(;(F:-<D,F2Kf<Xe6g,&
-<H,S10B3=M8Y^&-U:BbB[&cgD</#_:PR/[_aM:.a@e_f\e;#6-4?1O3.f:b=:=@
/LJRg1Rd)/5><AYJCX+HNeS#<]@AI[f^@+>LfDC87DJg3:gL17RIK<BN:RaRGgZ\
A3X@fb(X&Z3-+X8ZAg1\(FM+a.JJ(\7NOLa5A.))_aJCdZMCL_B3Y:0G#2M\<L?N
>@&KMU(>aL&:96W,]e4+#W+\CTC8F.>cS7aLae21>YR,N0/1,e;TT(?0@@>HFLS/
>aFBc)YLLU.NK9ACR/^0UQI^d^De:Hg]LM-_IL,MNcJLL,HVg4>cA^^08&_O?Id:
be:ISS,;A:d#;ZVXaI.NZd+^G/_&CJ;N37G_fNYX-31<^aGZ2T@D/bCW=2#DTKL3
IdE,Y;?:?IfOfHFYCGQ(](g0TFTYQD/25dRD+Y9e5V876N6eB.#7@H)H[^OW+<#+
10(Y1_a=\e[D?cCb2_\?>NY)FGL3O:35=B@FIZ+gLJ(6#A@D)^,6SD4GPKZRUTP#
6&4(FB,WgF:4JCGTPKCXQQ<Q)\6IGZ=F0HCF/dNP,1T&/Ha.C<#g&2N9#J9?<A<S
QYf#=N0?C\9Mc^?VR^d.1P_\]][L6.S+=ELG@+A=)@^@N;HLJ?R/9B1]]]6I]LKP
:5/.XeXP#4d>=8bBS=Y8YS3OQ50772d49ZK[7/IE\I,8]ZT:PE:fU8O22AY>314L
ac/cN6R5YQ[N_U=(&(\,ET3JVW?-5[d/a-)C@???0F&#1IFYe1.V--J;;c[NXX0a
f7[a(QC+M#d[U&Y?ZKdCQ7UV[SXRVfK,MR&?OK>^FP;M.fH7V0,.?X_e7HX@;+Z>
&G0V/3P-FR+_K4:fA>T]fF-NPFTWK&/^gA1gOGEUL7-Z2IG)P1K8C.>B?5Q<Fc_1
4T8_[=_Q0fcS1WXZ)Ra;_F3g-^aJ_F3>Ma\OCdf6UA;&ES_((;U3X[X80Og8W<4>
DZ:=:_T5<>,g92(0bFc2A8D&@cRTT4+b0-N,S)&e<,5/<gH+.C11G86Sd]Y<,_B@
]N8^b-#ZZPaB15[KTUe8eMG/,3X],4C;Aa[TgTIOb6c?HO_<MCM<00^MH:I=\gT(
O&=9cKICQ13CB[5]&W3,d?5,I.(.G]/((+Zd5[g4<@5=?]CVb@O3HSG\H6Y5#;]^
T=e/f9b>N/aI3eJ(N90PZ4D8;OVCYC=;]Y87(H?D?+8W3)3/c/3<X+BU[RQ18W\T
G[?C;H=N<-0NC.DSAP?PMURZ:<81+@)f<AQD_M24<&@6-_CW-8)9G[a,>,I/0M9)
S:g0:]1]@@J7^(/(QVI,Yd&Z8S=<D/S6B(FX?(M,F^I;?GGTdN/Q4K;d[26f&M/,
#G=P&XIF+HJM4&C@c;^9;7F:R8ZOU=Y^gL\#Ra6LbQ<TUM_M9=N69K^>e^(4\#1+
;1PNP&bY=+24US1004E;US6N^RcI8\SNJN/8:?GR6IY](\9UbbaRgV.fcS,3O5g\
BW(a5TKW89gO3bHQ10-LKSW_[Q7(#0+IQ,N38]Da#Y1,^>9Gb#/#]N4T)6L:38(M
A_G4g&1QO<.b8J75W/Ta[7:I_[_)#&U@_<Y5AR]dFT#8_E9AaFf1]NJ+CP\:3#\b
SbHF;8POBT.Y4SgM/c4UZCCYGA\.N[EPJMR;CFaYV&YYS-V2d-XbS?5MKJ1cd5bb
;9BLKcXP;11]VKB(ERcY)-G8UHE+A5SC4WC=R5bNfE/;5d8:0]FB&K@W-f?gZb#S
VZ3SSEddg0&KgYg_93(#=(=_.^,Rc-Q0;gfb/45U;XHc/2>Z5+<N1MOL_e&,1O0K
/5d?Ec1LQ^O,MXA(&)5XJH(O[BQYV/Y2c7T+<47VTKJ;[0?]-2g@,Z_UQ(YJQNGT
0U[46]4dIN88NUND[af?a^]&2EYRBY[;NONEO)66fa8(VUBSVMAdgY7/W[BIYdC8
R=E[R>SXIe[O2)(;;],8Y_M_72a_9\cBcG;b8+^cH<A^+D[7gT-/)Ge2ZXbC3/)L
3dB-\G=/#8P5FXX5?c42(bM@G-Ud&7\8d:f,P#QfQe6Dc8P@F_eBe.JS#Bg;f@W(
9ZN&V6?LSXMOb#cG]R8B#\QGe7PO-^MMIKe)C?42S+fD8)8dY+Be#+:DR7QVCCT/
D\4V4G)=]1#TXK/QIPL97\URdVEN6dZT?R<_@26>a>d3VfAb;GUbZf(Vf16]#MMf
bW&>K<45bQLBUE-H5/CP=:.C4SdOfI>5N>INSU1ZP>-^f?QDZ5^Z\F8157LR71eO
e=&L+-&>0/DUFNEK3/BEfJVZ\AWN+USgT+GGN16MXMOS35H1)22T]_dG^QA(bdC]
][_Z9]]6/KDQ#QbUa.Q&=Q>T+9IT0,V&J:3SLM6/>,]CZW[U=cG8?8K]XS;NKbEV
9_e.,bUYMM.0P93K/EB03B[6eW1gSOeZ-)3aZMDD(Vb9a@=49DeINOO\>ePc0E5Z
]D\^Y^CJF:0A82_VK;.O84C=U+6<NWXAY#=2PD12+P6]cD81,?3O>f+GfI7Sb([U
&;PWYTea+J^VOLI3[(+8_<&ODT8+g.L<ZKMVXK]66aY5D=;Q8<LI>WN[N#0<J9+2
A6;6J6&2IS@Q.TE)f^M3cTdC;>&Ed;:()+X\;4SV@,9R&:&c>H;/V#(4VEUQKEX\
;2^PA-c3dOeWL9c-8?M6H_:Md8UY;B5:JAg=JY>0Q,4,\MM@+;U+[3IFP7+FSbYZ
X+.)K4gH,S<CefJ@0#N2b,:-BHT7+>?=f#X+G)TQ1Z,QC3eR>VU4:?\ZPRXGK;O4
8;T?/c26I2Ke1:X&])-_BS\KSF-&TI[#]&@W7C[;N8C//@.J4/N(1YaE[^P&YICe
&)Mb#?a#NF-BE<YaWa/9deBCX[NeB64,,C-RFee\K^MeFJV#e[eH/HUS\PP.=ZBK
Ge&FYEE/CHEA465gV(@G38_:7E)YAR(M81DgF>D[D^GA@D(U/V;;eL^A3&NKZ#Q1
@g+;eV0FFWC=PH?&7.?fZ)>3NDN2^7a#M#:I@g19[[&+eF(8]Zb-b)D@G60dP\T6
+?.\<,\-UPNGLe\MeV]T@X[_,5I,@TM?B2I_]aV2#^BJM-/1(O,HY)HdZI2(=AJC
:_PQF9GT00bNDV6_C\.K\eE3bN</L;P?JZU[cBE2M^R109YQFY/&CYZ>I0R4V;.Y
dW69EfZ_=/DX]aML75C8@eC7(>O2XDfcL8U->R53V;9gWC//UN68@dcaB58DNA]7
3KCT.G;CH7&RW)JgGe@Z4f6cQ^>GNLbAY_QLC6D]KVF_+]a+VG#fBQ,c@\Z[]N2#
TK1_-OCQVa3WNXe9E(4EV(Y0GAR-B+N2=P56Q;.HeIL+e)1)9\<L(.-WL>7&#?QQ
Lf21g+(eD4#ULaAfSBS2Kg:Ud95:B/0T?d>bbJ.6U(J)?>N4RH4=c185\SB:^@7X
9M\gfKe>EJa(R(^?Fff&B(3AL]5M88-[Q(T^a+9@+6Ycb\]3SIC<aN/Ad25,+Z?b
2J0H_d[@H3.>AeT#2e^TJRV]ITV3NBM-e99\V=K&7E#A]5@YCWY>:DcM/[+LdUa.
P-@[gLB5]:OGMGB;#bJdSS>X2H#5ab[a.25E92dXJQRbD5G2]ff=D<)<F6W4_43Q
fGH7FHd;\6/AcNKF8fTGL?Z6MYXf=H?fZMg,Z1NA0G]]ZXb(9YUTb+@=E13K;gI@
T7cU<f0:43;@KC2)4YC1=LMAZKZNA?eg]RV+b=>^G7)Q?b#d_Cd]6YJ3DS#X9G59
EIG_5gKeYPQ9&Xce]HYZ&Wd19Z/N6?9?1g7NbMd2>R_)DH#a:RV+G^+<[YRBHY(I
(_H=>LDQ4RNED)g?G+e/5[0#I\7C)/T+0G-RbXF#(d2H\PQW9+VH7_>(XH;N7A:Y
MIe8(4HgV1?EcV=<@MA-H2(Bf]P?#H^Q2@GN?Td\EA3#:1cVJ@67^4eZ-P?[-QO=
Y6<6=9/Y96&c2.#M)S,S>00#TDDCN+(FPVZ(T#G?/L4)bP;eB/??.]OeOe(g<</\
&e64X^fWCR6)Z[I\W&6M7PTG9O9Q#D[&?Z2f6B3VLa3-PTF)#3VAS9b9&?6(e\5\
QWAPM8439ACA.\^dH=g0_OC3G@X=2gF7eNR(6C:+O=\65g-:]ZM^b+I?2bgT:0-K
Qc>P8c,SMEb6:S<;K7_93A\8.@d:JQa0R.@eGSBQEFE2O6]]=;W#b-;4IXc,8C:G
=DHU@M+T(TZc6_B.1?+[R.<^AX;Cc.aAD66LRH,eY+N<E1Z@c\BO5[aGOIMe5]Bb
^fG@,=A_=L(5,:0.VWD7fNgdd(MS4N99]M[fGdP52NJ]HMJd<SVB5g5W?3T)2egI
db38T@dBE-Z;HXeD^_/&AG:<[Q]3+UMbQGWIG:GA>:19O&)<^/B+<G7&S.AOOF=V
F0ceSRFb0-VGZI(Y8V2<Y=cK[gQX6Y<5897+W[@+9L>BSG>Q5B07IcbBa[J#\)7?
a\&)J)\,.Ac?+C(+Q,I?(bKP.]eG8N2\GJe0\\a/0cWPg.K-),#[]\2)U._1_RSC
2+JLH2SV;&[.^+gfAU3Ub\cJ,ZCTdGU?:e78HU0P]YLPDB?V[\/I<JA7IS3=1(R&
&P72?gX,(UX;3E8QW<,,K[]JK>M29d=L[^QR&a[8F;CLM/E1RfL&<ac,QHT;Na^a
KOgdB-XU8fT#@)PN0PBN;<TZ2cY&3HC?^QU>^&P;P_R-HY1J,T:_AZD)@DA\R<5=
a2a]UYT^fae:g]ee<8=gKbDf)eF5eb7\Z=(QIXAf;D[fA4,O1&6JPI&R5UX,Y[,?
F@M:\F31[EDd;M,:Yb&@.[[]3&b+W/1A61c>ZA:,<]1/S^JDT4IPOb7=\ZKQAQ52
D5T;&cD=VAXQaC_RAGd-EC_@-VXFDbcXGZbV[<FgL_XC;a.R&V)11B70/BgfTE=?
DgG2@WUg&8S8IWM[MHY@5O4)2?FH[Kb@1D[=b02FKcePSfGUX.NRcgH_@dF8E?#9
gH4Z9\YfFHRKH2D9FX@fCHf.S)<Rc^_SS^FDA=aV\:C@=;T>X2eNWc.:[CEP\/b^
8@-]WI_D3-^D855O@#Y,IOc,F#DNO/QD?<M4ef)<b>ADTP#_(E#MC_eFW&<)CHG+
,:e&JE-/PfLOBbb-ZFF#)_^KU6^FWC8U\6,B.,YbKI/;X[27FCDUVcKH:38FRS-I
A:4AH&(8E7R<2?^_E.gC;P)ID0+LV4B5:L[&D:dGcP\RBNX,D0>OaEJaf;;UZN9^
;TCMIZW-4fM581H>6J)<CHeYSASAP7./>I@6Sc(?[(d;\/<8-8]OQ<?-I#IL:<).
UO\L/O^=eMD;]2d;-XDI#4#KIg;fX72dN3WcMVC[eeN/6O^X]<+b<D.<W[d];IJ:
B;J4Q@&fgKefCbCOQ28C.#3-[QW@Vf,9CCJIDRE/HM-:&3DH@aeYV?cG-d+e(L94
b=X-[^f6),^H2RAb8LTHSVO6>]0Q2O)]7_8+DCeWc5CZM0UOa&H8fR=6@+KD#8=&
.)T#2]A_H[>M+NbM?2TAFM@-(09O(>;QJ=gW/aa-3_?)XAXX-Z5J)9^IYZWC,X_d
?XOUGWe15,MUK32X+M8.GGfc;ODagccPbP7e)[1^RU[HQA(W0)RG@4M=5faAU9_K
CA9I]&(SDD[SY?<c,dg7@8HgI:ZNHZ1fC]T88+;.@V6.=&0V&Q-gaI<<HJe?=#:5
9X>D43.(P^bTKDJ2g5,b=,4Xc()3&_c7SL1a;^eGf+1RZcZV_QA4-V+0NaN/E6La
@Ue/V4W==XPKJH,,bUC=T/__R2=>HHgA2LA>(G(Z,fQ^.#GM/\f-C+RG&eI9Fa/C
FeB(^T&).]<A0aATV(^;ScN.OY6:[/<WL<D?AbeN48c^HRc2aab2U@Z64:\b1BH4
P/cVbR;G<a((8N2OZ?L3@L<e27JbF+2O9H3@B?-IHE1DdUf/40c]fBB0A&WcRIBM
>LI_1dYZR]g90@3BW&:C<D\3-78UScM^3fH#9W_?CI)D:HBKga)e]/@DRRfJT0/d
Nb(>a/MKHXOXc>:N]a@K@?X9ED504?QIHH=EHTIY1(,>RN/4R#.]IZ2N[Y&EU>/<
Q8B^+#C;/E^L0_5f.X+gZ+#>bJbdPE-)7=VMGIC49Ve>->]D[XHFR;S?<&-HGVBd
9C0aC)aD5>e]CS4X_Z[(a4b+f?4U697TELgH36NJ25^>2E]@PP&)+L/R).,V0CJ-
Q&VLeAR;#)P6T0IM4aH=^32.<CY2;VLH.]Z=Hb1L_=-_=bUH3Vb.R>gDH,#B==S\
TCf:AI.e&)+?PI(SRAC=5YG0P_H-44.D8WJfMJgE+O_/P7If87DGHT4@g##B/^IH
5-cLO:EQMGAG70fEgL>9=M-eQKGMYPU[=7]f+WE-L8J>IbI1A1)P3J#-^5b[c)eH
=2[9ILK?Z/CHKN)fK8cdb8gaN?9c3S>7Id,<ZN@=6>U=CdLXKU/YVUc.<SAKd.FW
=X_2aIH<XW>S/6YH14XWd\-d[CY(,9abgL(23Z]YCJ\@Ca]Sc2EK:69LK5^PTHR=
IO)4DAX>^297C?EHaE-BQ1OETZ43+=dPTMPZZ2JJ;,e:>=XfgJag_+H8._\X(>/<
R)QW&DQNNG7EH>VX[+1L.-PP(6/3JI[:.)K>\-EZS(<cEfP_T-&:F9,a,D(dTYd.
1RSQ[/2:6(P2/@@9547NF_2X/NYI:JZ9_3CLbMGQ=<Y]UNRZUR]7f)[C>^1,c&8=
(@RTERNF,ISbP4<@D7A844dbRcJW<\&@UYe)dI>?cVSL)([UU^1RY67)-]1K2b^d
GPVP\gGGL<@He8=HCF[+=<VeL.W43VEZ83,/-Zg[)[3<A)EQ_(ec3[CX>/-0NQI6
H[7RdG_[[U\;>f<ML>IJQ;)c9I#f45S;,;XNM+GLX+I3^P@=&c>L[^/J0+OHE/\G
Ta_A+KE0A8[BeX<\:PZ/_=g(>gJ=-)I\E9YZ.3&DF>&]6BEBDZK^=(EKVM_:=9=D
H]OJQ@1N_1H<X)gS?5V?V\57X/2N/79dT<?Nc)3JONGRf/U)V2O:@=7QDFf6:g8-
:(QF+&c8H:7TB0KB]J_D;H<_VM2\@K=&V#7JSN1bg](>:[BP1KYRCdV:gJ0>AR#B
EQeJ8NIRL);(>Q@@-+V;FZ5.EMc98>44Qa/Y>f.,^(bIE0(U>C4#>&/ceL&2WgZC
=>[L_R4K[Y5IY4#a\/XH^)Z[4,&Gbe0^7N&7eR2<M-96@U-K9VT=5MLfJ].6#P=I
,<0Z1?]JFR)=_\0K;5;1H^Q2^a(d0Af]+3(3_\eK8UHJP;;R+JbW[\G-/1QAEBCA
acO(\EL(#U^:<TPd83B=.5gJbbBM?cIF:K^dZO&O:f3eG\/LXD#M>LTdBI]_@Ab2
VQ;e@e1:/=AL4(-7#de-Zb3G4^X-K<5\P#NdBU]GG>PVQU#S@BbXN;<GUe5:8?](
>)BHD9YL8].=IK4>-EOQP73-;?]eQJ5D,g>f(-bX&U/+\H2&C.7#);/(JBc(QE.>
g_,1<>BC=__4Adb9?_-34T_dB-B#,M2+L=]CL2@3]1]9CaE0P-@[D7ATB;[/Qd4N
^c9aWG(-IQ9gH(B0#AP:.2PE=HaXe0^&MBC_;PG3\U,#^F-)5<ZE#[O7Hf\KBc9W
\;+-G8Ye.F\f.f@Na\@UCW=K=P&&f/PBYOJ1NBI[b34]?3K0ON<YbaFY+<->4/S1
UL?S6G8P/><\cbV_6Kg7DYWWM)L5TOC4O@OAg33P/5#\^8B6f9dAJbf8UCUQ=\[F
4Qg1FZdGAPg<ZTGgI8EU<EJWSN2S&[(S:c_U]\ME7]_QPVNC[Z7@=WWP;02+fFRX
()f1AK8,D7D2KAE_U5.D91dI>B_AK<a7,Z1GQ7F9]^>JNQAXN1XHAcT5VE+4a(.d
#N2XSQ53>H,@?AL#.3\>\R5BVYG278?&04+0V^^6f@a&.JfcS=WOY)1=aHab1T[;
TAF)6^6;8WgLSe@2/\07VRALa:@IW5K?L+_0?3[Vd?MGL^P&g&7d1-G7B/K>\/9L
<bg,8F/2PJD&M6RQ@@/NL>8LAW7a?0e\F\;]BU<&^W7BP@Pg>IW6[(F[SaDOG3NQ
&F61V\GcgJ>a8]C]6[-DL+\@3@PI2dF_NZ8+LMT+WYM=5U)TZ-YKR/4V75O1DXX^
])d+5I=a.]YM:O)11GfKL)B,VW;gEU&F\6)73/c?bH]XFOX\]=SHd@+a[]Wgb3f)
U2?e>YdQ4HP)>^gL,F702Ke0]ZedM_b=W@\_IFQB?YDH)L@;>d\&97IFYSV5cQDe
EU.+P>R0-C.aK<>+&JR1_BY^I,VT=FI0>Y&/d7@IK-Y(LJ).NCf2ECUCJZFfU3N<
_N\3GG-97R(.d&C8aC.?E<\G[JL\JC0#/LE\d2cCfQ^5T-O,d^_[]#J)AAHF5@M\
+OE^W(N_K>@6ADCK)#PDBJ1NG8@Z7Z_BZPNT0:MU?RBb/=F?76+Cc452T?1@XgDd
)eFe8bTN_60K3a:]P@LLYE+<<AgUM@7V&gX)I#BKQXBF,WBA]6_SJ&f@FgGB.5WL
HGS75)I?S=Og4]MBaIeD(46G+b@,J<VfI^S)S-c6?aBIg&-0;\T7FKW0e^0I4b\]
5d9XJb+&cA0MHdM3(>33TPH>O#9T8GP=2)]K40J)F,T6,Yc(caIRAKDF;6PK5#.#
TBAOV?/K[e1>^>S_B&UJC(706;VU_-UPNKXUeKfT_J(1-)]G<T6P[?1UHb0]1gX.
<C&1:NQ-^N^?>EC[^M9;YHJ5=Ye#JRUd,+4Ke-T[Q4.gK6G;/Be0H;;W?CL[cMg_
[XDcSSN\Ha]U3bI11_(]Db@Q0;Z=Y^G30/2?:d(aE.EK2,Of2D_1K=7)U)5BeGTE
R-,;6MRL#E(@LI_:Rd@]SQC:LQ:NN.\f-F)Y1H/VC_#(Ge9(=9>@@3565,)XN_Y0
aR7E@ZWQ]7]+d:NGW6I;._I>Q+FDBINWFVA(Y5[5S7-9R^>P.;Ye^07-M(V:V+aG
BAe)FD.2EF7S3SdJ[X/T)Da.563#L;B7fa3D]JH=/5fGB1[&\N2C;>3WNKOX/RDV
U5/8MZM+eF0/ZQ1)H@gV_OJ:BYc)#=EPCIS0>.2.P04)2)PM#IW_EaND9eA>ONL2
-KbX,HBfUdVL779T2,,94aS;/1HQRQg96W?(eE7.8a1Md^eH]3>JOMdD^5>^ZT/?
&_<3B4F@41=c1D-/;3<a8Of5K7RXg>;de?\IJVd9D@2H]e[I^HKA6\A_[7K,+_R/
WK@GJ5.OOJ+A3UU:AXZ.&Yc3>G+PYM?NLW3\V>TVKLYE_L:N?C0;La4AS;N5LX+:
5^W_fJ?6?0bX80\AJY8e:+M<LK[Y8_5W[-1:Y(Z:=\V5b/CFRW#MU?I-(W6f6Kd8
).[=4(R0BME0ME/>DX7D5)91]C(8XWc>Y[f^ZLI(6P.)8=)dMLIOK:-5.9&G2eg(
Y</#ZDb604(+OS#K\[7_BfX./ce3DM?#XKYFW9VHPZ9?(N-I8]cJ\&6=c>T@g[NJ
(eF/?[DPNQFE:eK0:Z=D;]@=LHCbg7,VAVb\2YI<T_6D?e7[<(1=7O==3&PU.JFP
S_+7IX)#&J()8^\-VFZU0R8dTSd]^LR3GRY+)?Y.geA@SZR##_V69]@gYU8-+@g=
^N)&\L8-\Y5<JD9:Lf176FMG/]Pa9g@VXf?;7W;Y1]b+Q2><g8P\89V<7)c#Q/PK
dfR8&_fVacV[@#XV5edF>KV73WLJEIW^9_9=NXPR[75aO:^J@3T>/g-QGSH\F4(6
(+1cW-].HYX3\J.QL;a>0M##VZGGN#_SWH9,Ne:cO;9UaA:EK.7MG?]KC=4Yb3e)
?>bTd_H.I]AN,([#eJ^JTTe9dF^:6I2UJ=Z][7.(B07T(TZ>SgJB1Qb7R8Qc[QQW
;^6.K=&Q.>_IJN(-;10()O.d26]:]_6^e-8(,U4T^,Q1D42FP1ATR1fF>E?D(VZN
JPV\C]]]fE;U87A+V:<E@K\II3NW7IPYb+-MKB@3QH[0d@F1B7)-3\:_MbRFgBdY
YE9f.R[.a=W02TY59Ce;I,/@,Vg#S4@.bX_>(cU8R;Ia3@>[Wg<AM=K\NbJXdZ(,
1c/LR\QfBP\=T]<O9EU1^&?#[(YSAM+>[Dd-03/C6NYO_F0<8+YVW8OL^0=Db]eK
KIOQG,M:(-//XP&A&4AQ/:@(KcdB<4aSX+Ia86e/:^[K8I-R+[gfWZ6EYBPHDVVa
XX\aEc#cb^?I;9c<8W@\4d&?GL1_E;&Y=<Y]@MR)G)G40b66_:Bc1)I:7M;5(+d3
L?-KF]-5-VDE71?W65_NeXIfD>6ABD4R2c&N^4D^SfdH]UAW<HT-@0A;5ZdM0=2P
V=[^/Y1eXE]egf8+I22ZfJH_7U2HIcL[:LVD1f<VM.T?G86cTZ_aPDZC67[\^a<.
9D.4H5a9Zg<1YG?=BV@3/@_cd(52KVDP,=4eW_HPb#/=8Dcd[SQK?&,WBeN/4>7[
8QV60W_b8V2+?3E7bN:76P<dW[FJWKT0E8?P#;MXHcfMc@:Wf=BIDL@7-3IgAK4^
D50c@DH[.@K#W^_>R_J@ZHQM^/O_NQCLf2=RR5g8PBKPcDN[C<bbL?5Zc4<-=Db(
Ff7L/-U@e[ge8J7)]gSEeU;.OKGD6LRO8)ETL]-/SLQC6[U/@Y37c>BY50f[cI52
V3CJTHS4#(Eb/eCY,+V3_.a8YbNFXQOZ_P65QF>gI9]cKga1=,QU-&O.I8BG0+[E
P8a7.6W+cCC?D.^I27KfUD:2RUfFMKNE.D&#FCYM_&dH(b4UKT?RK9VNbf7E7E]E
CgMV&^^BG@4Da(F.cQ/UHaMaY</<.K8Sg_^/GYLe3QJ#MB5MJ/0[O;+Y@2NQG.Sa
?N-6CSaYEN/^V9.dH>5\;[97gISC^f0-L/5)\Ng?a_O=WV,If.<[TgTPMD8S0P+/
#QVT1I&70#L-V/F=6;e:RA2],KGF,X64T//+(IbQf5]F+A3SW@76AY\_#c?E:?8c
3T++JK1]\0=CgDUaBbF[<M;;f\?L@d3BN)W+bQI#)(_C,Cg1QfA??_/+JG]V;3B8
a,3J^ecJ-C\@/YZggQD<X;(4N0A^1[:fU>?B0dXE\4@D5/JP((cNZ0Ic):IJTID9
UZCIK.T+H9aa.Y7@Ie8PRM[KQ<P6PHLSBL+?1YC3Pe5R:Rf:#O\VOLKO__C5PGbb
8AbT;V.QgSLWI\?N.W:IA6E(2)U&b?G57V_9H=5W=)7S,N\3\G<U_>,(#@+VfIYb
U/3R#<+#gUQgF+:c=^V8A#/;B<=HCSG:0g4^^,LHLQH_N[Y446HMF.T)>#eN&HQQ
A-;g:<.>LM&Q8N<[N77ACK?L.+;Xe@b<1[[ZaO7ag]SB5)fa>Q9a?&)MHX)4^&eF
24Sg;\g[UAU?@g06=?V[7Y8A4@-aeL@]CA5:^.(SIe8[=2(b6S11O)T53K..:FMb
3X<#I0cPM4BHEETRb1\)\<<7<=/V]P(W^-Q_K/KZT(dF4)E0bbO-4@4S)TS?\&=:
3fNJYX)F(?eCI+U,N,K#.^FGMC>QfL1aN_=C:I<Gb?dg:<&1&<_0Cf=3HM2RXT=6
Dg(;V[T0NKJ181aTXQ3<0K<\CABbLa?1<XN\dKaP&\.[MY&NY_.b:(U&)7[1SM5.
B:]b9UId@.Q(Pf]Q]SG,;21e+&P&^g:I.ZSYgZ0)(00J9H0#ZV/Dc[_A2Sd:-?WC
NIMF4<2OH^/;NYX8KS[9&eJS0??/VD)36XF.O(f?^B(PVZ-gB^0a_C@H;.KA\+ZJ
.B\4eOZG,V2D1X\>T/U6:Jg)PZV\/\QcKgR?YE35/Y56RZU<YBL]\7P6U<1^G[EL
X1-WO/4.O#EH1M:(Y^-8Xa=cDJDGLCe3gbI7cGPCJ>XTUXbZ/[f^Z8.&5R3Yf9:<
@\<0XD,2GaNA#1QPG43#3DGAD4;W#WZ.ZLfdV3_bccEBB(//SB]3^9F;T<MG-TbR
G6SBIPgTJ&/aJ=DA?#5BS@(GOG@UIgAX)e0Cc.Ya=5(/_ZHT(#CVJYT?6);\3\D\
Va+bY><-bBJ@,-SgF7)BVG0J(5,bLOD<18(?]ZFO0&OPSc6)7IP<523eI]a94Ec7
169V(N7Z\EPR)0ZE[++\PHS\3a4Z;d[.]^P&d[f78>^V(3R[[0L)K+T44>>WH@@L
<7f_@C/3X]@[1=IQKMF>Y6V9P4V#AN9W_cWQ^/J@dZ[^e+7)OgF\34ZJE.gD>BFQ
a/[QE8,3TO5T?GENF^B\Q\I-1(/JGO=]Z=Va(LaFUC1I2P:.6<^?);\XdXeNb3We
C3MMb[WL\CLc+=K,VZ:KF355.E[L\0WTOJ77ZIFZO,O/C]]F__SRgD9:bBBA7T#;
22?,J<FP7TfgI[M+5F&G)ZG7BWBbC7NK&,e>\gR/e+L\JJ/DB@061\)ZL0;b,H5V
N_0d:LLZ^-R+1Y2(bV[SQ\gPHINVX4T16-<;-/d7f]3gVI=SW05DAIBG^M)XM5PP
PAgFb,GP-^XKTOg8V64\_a<;DD\H\TG.,Xb7;QK7=R4LNa;X(X,AXT5IaO)C:4Rd
Bg2G(3]XO1JU10ccI,OO9:_;H52f9EK<#.EP-1S;>Y?MGC&:;bcb;H(eT]/g?2UJ
/P2_d3Uf0D-WVC[G35K1.ReYf7VB+aE13aI(,A0OYI2B66a-UUHK+a]?Q]D;Tb>D
0EAWeFTU\O<X]g72bUEIFe^#IK]G,8+X\R-D(0MS=9.#&@^PP6Q2[VPZgV+V30>;
6X_MHPWX,,5(a,V6b_/^\5B::CLK41ZR[H2.::(M(^W24#47W;VR(LZ-69.QLe9(
ZK>6QI3bRM8LV^4Zg[2T4P0I4]^&Dg8/?G6S\2)76SI@CF2bQa5Ic/I[FE/H^_Y9
SY026CgB+AH174K9-9N)1\E^WEGN0>RO.X8/]Vg[+<252Xg_K[Q+I9)J-?-_L2]R
H_<XH(:LZ;H:WLOI(_Q&CZ-T>cTc5O3NX^31FBODcX-A]8[2d,S/Z7<<B62+d<DH
4=,A><,119#H.=8bJ=S0+(4)&ef-c)([)7a=,]fCC>OC^K2UMA5I5@004,;>+/a4
<,c=71N,@a8B;W[&2VJ-#DLAM8N\O-XR[2T#>+JXQ+N.NE:N.;GA\aLb\ZB)Xa5e
e?[4a3,JJHCE05^AS_)7>-(KGfGd,Y&gZ);g(VWT3GQ\4F8JG8,[S^Vg[YK?COeQ
-H0^bPB)#B-7)ZNAL9<>-G\7:G3YJe_Y^KN@>V(6\6>I3U.2RAgB.-:78@Q9Sb]e
UFZ^cfa2]U4<8^8IaA(E1]N4K/[/b-@5-(_TB?25<L<a7BOf):.Q+E&H:gAgP,R&
1_+8BN;;3/[9KU^3cQ9cXE30d-&N5NW1X);M-4H,MALf3(\VS5F@]a.0H21e\DO6
<[1P.2HJFKa27g.bRFQ#IAL:4S+[(RQHF)0<gAf\:I,Y-6(A1)@&@@ga-=V>be<U
WHPd5bWQXJcS)?0BO_2XE>TWM\P^TEFe(0+,R6c^:6).(]PGSa@M-XC=dd(0HL,Q
f;NAOISIC..&RAc;)R<YLYAd:H7NQY_^dK<=?(;E=,K/UBe1PJ.F<8adW)A8eH&R
gPM^Fa(DIFXg=D/_YP:bb?GaF[O+T&(-TP^9O2#;AXMg\RNeNP8F?UdK58T5JDWF
cOF1ZFWW@aON(MS(/P.#W7M:gGL-gI>1_)a]<5R7g6d:VWLV6dDgd<<e+0cOX68A
P<J84[&73KKI;2Y]^QP;_BfPGNHN#D8A<S[:08bcJ/YNZ1P)GY=M;gQ9\TP2]Qe7
)c)DVZ#4@QdZd=L9=eXdbKNb[P/ZfT0a?c05&=D:BW-B?,+[?;0_;c:&L_0A>#4g
FMAZfL-LC60IZQDF:T]QO1aFQXgC,YGdcPMS>6aKN+>WadG965O@/5VID)W9E#^W
7B8R5-aM\Q7&Q5&f;,C=5V6P;b\K+C[OK_OC(\M>Ca?9()8RY=3gf2b[<dBU8B-Y
I=(@0GdCX:_7-gRe1.e4G]FY9@K20MDGTZ#OR>c)IOA\.#gW:eOSFPc/5WDX>HF)
F2;_OUAXU7BZDRa)(X+3Z7W@\I,b=b@)GRG?PWc_dCP0[Q?XED9NIaH[;=@LQ?J_
^8=RP^3gB#)Z]b5bd^\C3cJ-fCb3+GW.Yc5g^E8Ta]CG^;<@eMHMOFG9=53)][Pc
ZNV==MQMcIOKHEJ(H;^P[c_VD+1N4MTb;acH9V-ZXWZ[fB+:XdGDd1EZ/e3(L^<X
MTHHPVQTV2L@OZB+.JU+Ib++0dXC2@W_OA[>\gCMaQI9>g1-M<F\79bc@\0IXBXA
29A@&SP.XL;E3dgQGb]S9Y[Q3406XPZJNGK+A3);DRHPO:5),1CbfLY37(/L)V,P
d(WZgBW2c>]5UP_\V?,K=8LKW@a,)G[<\1D;H1.f4^X,RKJ9K5-A(9\9E=)RW^Xe
>2JM#7WLe^+\.a/PAc9;fWPQ,0#EKT[I0H>W>gfZ0R:?C28_<Nc;P3#5g(4-9F17
f^>3E&QXA?JU#^]^V/#3PgKU=N.Ic_#@@Q@2R;-<#)S0868&&<=2S5g^cbVR]87+
YHc=;e4:I#A#.M]AVQ^;XaO[]MUI(>DRB0TbQTU,_W7U3RF=50=YW+DW6U^AK3BQ
M>2)CS^>cc6EFD2MdF1>SV(LUX#QHC[MXe>NBQY=PGd=\V-f,F8S\QY2a=;<^ZF3
0c?S)X^Q\AJQ2?VVXA]3g9]Q8C0,)4XD?(<S=RVfC_#6LQ07cDC^XGTL</:/(C4-
dC]KSNRbU9Ie&K&H76GE-d2N]=+3-:.917L,fSNS^JRXaUOF,F].NSZ<RL^[-]VJ
dPMLT+OHV3JHN2V(EE>2c@>TN\U?4PK+Y+#2BY<S^a48,O8+O?SdF\NC6],9CgJP
KN6FS-.:-HJ:=>\:Z<UD&N:=GYF8_=Y]197&MOF8Ia@0gG9FUOX/Vd8;6K&24LR&
D,:Z#gTY)W9f[9ed03CP/D.S]3G4B?8-2FG,/U&XLCdbZdBb,)+&WID=C>E(S4R+
>8S3>Kg.2b[Z,;D@feb^9SWCANR1D;@2\;^bdbg#1G)K_Sf(U[H,7LNX9:e4aca>
^)=N#<P/ISW7&>/4&(Ed1gcU9)5,LKIX+3F<g-a++8<UIB9EZfcOg;d]4UN7LNN@
AO]dAH;8P4UWfWR9_P;QMgWM@Ic]-#/]N5J.OHKgHCae1](-;5QI;bR+XT/AQ2C(
-eY5&fXE@@@cS9@Q([7;:CI+XH[RS]a^L-g#GVH-4V@-a59)Q=2A@]9).D2LAH5N
UD=2[8ZHXB+Y\;L7R+@a]8V]GeF>eeW59R+?M1C:a_:85Y.WaFbLEKXF[>aW@d/[
>D;Z,Ofg>W&:Ib,P+)4_##:[TT1M9>B.X#DDK7IdbKa9BY,E:Bg>Q[:Q&Dg#A\bA
B#>OM]G<T@GPaDZN.A>DbP958)3?Y4DRNXc5,Jg2C;d(X3,Q<M8ADDXR-Kd7<5;R
4bL5XR.T&>6W@/<H=bZS_,KJGYTNGgH[E?Z9TT[>9^RG)fV_MIXBA-^Ke[:\:deU
5&]>[a50J&aGL/dd73^@dZXSJ,N99_<6Q;aT.SbM^>280SU+:IBN\)LSH6OQ0J8Z
@:80L6(N(Me2BVV4abQ<69fSS0[M:_K<&^Fb9Zc:f]fD_Zd_ECN@OM+A:Y726GS5
^N(=G_]DOH84+=)SJMPXJ8)/a2A)6.,S,KM,I_I\A6-H&5CTQ8I.BE,HS^#IJZ-Z
3FYF?F1U9)XDR):WEFEa<A<\O8RPG+XJF]De07:7>ZHbbc=Tb+<eDe<YSKVQQ1MX
6](_JNf8WUggRFI.0)F>CVA[.BK0>89X<G@(VY/I1,a4]dWMG,W]@=0LCP.N;D>_
\KR3C;O9/T6g2B+8OcQ[_+UdJb\HRd0SP?.II;W/1BY4MM=T8UD&#)WM/O=5Mea;
FF(-@f=8-P6Y=&VU::Y)4@bc_GD6K8:2ZJ+UY6+)7/R<W7]Rc5c@Yce/fTgI\V5^
e]7&I5O+\fBba.VbQ^V:+Ve<GMf_2IY]Q-;1d5Fd+59Z^?LQSc:H67>=(1<@8a(R
0L#?QDL@0QLL]^?6@F)LSTH7AZ:L;K,[.ZH4J2UB17+)Rf/92c1J/,2QgEB.K;W[
VNGRNA6)=,8FB9G5VD(f#cIFX3TQ\V[;#7LX43Pbd=S^6#W7[S,O6V>@\6B1X/0V
.K>Tcb=Q6[,YL7Vf?6O-b,^=QQL37^eNAO>gXB2d8L6Zc2-QYF1H\d-dGSW+38)>
<.@[X;S4c3:/5O&Kf+NU]1WTb8>9K]&O2)9A>2.@4/+C@8X6HXF.cPM^<X54CI.[
X[-MPY7^6FYL\ITa05+)9J.fM75&GJ)5_+^0&bcGOXGPQ2Qg]4VC>)dU2LXAeb]7
4RSY?.\(R@feaP@P+CcV;#A:b)SLXSb(#]?1Z3=UMTG=NWe84D-[^eDCK)V&56;M
IOGX>7PI8HY8M8/]_HM9)@_.1M_((WT+#YM6W@RT#:4Wb?=[N:&8NW@7fAQM=_dW
B6DEcT.&GF#S5TUI2HdW]Z0V<QQ)M^H34#ab:;E]WeR,bH+e?CRVg?1V&a,V71?-
fO]XWNE58@dc?/>,9f_:/9JZ&f)12;_4N\KcUB;2+PDE2H](FF=#)<U6aB(6.J:L
=2>?V0#9CN@S14e_Kc(-ED;Ncc^^;41-9Ve@FcY?G:ef_Ja\Aee<\:IV)PUJ9>XP
DPc;:F8TEd<H2IN.[+;-83aB6H(ILd<X\;A@(G[Sb#KXPBd02D>dUBb2Xdf<INVO
C@e.VQ8US[E_9=b/8+EFUW0V-Y[&WOG2EXe-S5L^)O<Hf#>MTYFFH7;8eC7_/GI7
E:6OYe5MbJ2gI4bEG9@_AOVfZ=g?/#aIPab,Wd>QK#@LQ.OW06R-_@FD(f_JBAOg
9._RKT.^KO3Z^[Td_-#@<+T(e@=F(O0T@;SCLS4H>)EK-XTO6Z\IFgH=BTc9g1KZ
=[>NR(gZ2NS0NbA=Q,GBd3^UANJS)/(TZ@0,cJ+AU@I&?G,7N>Q<J49H,-a]AB9e
Z\D3a_Cb3]/eRX,>d@BAB#[,6_[804E<ED^3:IM_60GC&J;e^e(1E=6/IXY46F[L
<=HM-59d4-[>AFC2KCdD7+67ET+W)3\=1\fUTXWQI)FJ#XV\R9eXV^f#+1C8C)0C
E)M(T4DYZGMaY.\UKI\5NbE46UBO7CV]0,bFgVJVC5JHeN,VK&QgQ[Q12N5.8,3[
-_@U=5;Q(c3-W8MIG\YS?W]ARL0P5R-DQTOfg0L;Z74)O@2->+/6<3dJX([Re2L1
A=KSF-3=(KT,0EPAJJ&QRYYP@ZXUf_LDge>f@e/5Jb,3.VS-)=5/1TfDIe1H0XQ?
V5Y9KFaP_AAN_.EP9)#_AI93.URNV=G#YKXK9,E:EB<dbT6G9?;NU=JQe[TQ7DE@
QESdHD##-IA<G9S#dSQ>#J859;9b=22d94-&A8N\,M_faQ@NK?G]<#),N)b39J8;
9d@._^;V+-Y+NI.I^YW:\aD,(Z3YgSZ\H8@?8CUJ,F^.ZWPDTG3SZSc@IWA+6MZf
b)EV-WX@HK4WA^?+#LC3/XJ_#gN50OeDDG[UIMUFECWF^a@ILG>>XE;QBW60+X-)
(OC&J\CR1Y1H76R)C2[Z[H#48egDBCL_8HVIS4MF[+&B#@J)fR@MH0K(B08J3:7g
:HN(HHY0cALJMF4/I@:(RW8fS-<-J1OF43aLZJf:c/:-P0OOSO+\KI[G0R+;[16#
KP:^ZV3)Va-ENc-L8>VKU,#6Y6B&4ZIMgHeJR32dE-IP69=+(/:V9W#,X10.LH#c
LAb6RdaWZ8MACcV)D2DH]CMZ27:WB6>M@SEFGK4D9T0I(3WQ/\Ag<,ACQXHK)>G7
&0RAC)\be&gI83g&&fa8b)XXH2TI?6DPVc><I+.^+,/Z;(7=-Q9:;PW80+6\L>,S
e#X5=L#\0>:d<X:OeRdI?XfK(6#c>OCbCG-d50V^/)e[,:^eI/J]>:HO0>Hd9K>d
<U??feJ[_\IFG/f<C.K>VVHX=A>Q#QT5\@M;a&SQ6@((KYFOfI52.@^cYGRHZ5-O
3e0;+&4):bYd\_:N7,COCU#KYI14<Q0/d8\aGO[d_WR-,aG=bWXFCM7CH[c)e_0B
J+>S[\L#F\AAM?X(COM9R-NDE7/b(/>)C3OdTZ?cb7,?0MPF[NO;UM^,C+RK;[]S
_D@8A;S>dcF?.@[9OH?&.C\>e4R1.4;NER^9a46+gCNA74B]XdLPRQH3H-:WDZ(H
U(#cKAMCX>XCZ)TF+DWR+7GJa6c;2L/0L.=I4&N0??\>N9fA7AEg8D9.3M2J-)Qe
/2+eWH7X6OQc5P)cC&_1#@J&^[F<BM0BPB[ID.)a)@+<CZ1ab+XO,R4b)LfWG[Y_
IN3LC/[d;YLP?a-AM/gRO;#][>TGC4aM8H@3VaCE8PCYeD#C#;-?F+eEgYc;V<#I
AAZGV)DE#,_Q<5;<@^+4@[bLRBa7aLH].K_0QA@dN&/966&C9;9?KF(FE_QgJ>;(
4Ga;Pea.fI<1da[JYCA\\0aZ>eSPG;96gE)=6[ZPZ&QJTYBeW=)dV;([a/LS<H@L
[aZRE/]^9?)3\+X..UCYdAdf=H9F7(fXI@B]-738E;6\T2Mc9L,HKR^96]GgbeaN
SAaUJDV@3V8XdGbG,V@P.]@FeSfd+CVU]3a06-]&G-6^V8f>XHWg>fZP\R@;,LS5
N6V]C//UR@^Z:.0B<aYA0Zb4@L2E:cc65QfSaGeQd[fZU6352N)1&\2S[:dES(:?
a4f79&_MV5C>Vd&+G>]CYZ?2[)#]f.222,1HQ)(6Q2:T_?Z2BAT8:#PU[9=N1/bP
bc;W#^^\0bB9S?B+E3c6]gBE6ZeKB/02=PLA32^@NFY5&=O@Q?a&PX/f7M2;TQ+Y
>P\QaD/67N\BC),Q\9]=eCQ(FN7^(N8gb+3^@QV0POAVf?P0Z9:I,HRg,J6SA8ZX
=XG)4/?1>HgY^6K^^UZ8Q^VWN8W=M&5_Q+7;LE[#84QT;ZaUBb\HRe]@&<ZJAPBM
LUDZ7)baDQPX>CY?5A-OO=7e43/<8(7(1f[CATYTfg\(M;JW-,+IeKYI0C5A^efN
,/0@dRMCM7^SVJMRO5YERIA,(><]1bQ8?X1V8_D-/D+O@?&D_VFU:^D15fS?G7=5
R\bD[O/Z/(4F#?<K2P/5V5Dag3fSQ-WK9OE+fd\.B+XE@I-f5]AD1.&Eecb8.AU6
;g4[6Y=F1D-H3M5U=14+__L+H<?PJP5PWZ8<;U@g:b.3eYAN_YN;;-W#68KRJD40
K<f?YgC>age/Z<K;#VD2IX\e1XcgR_5g<ZKdNTc&LZG5OS0Xf,IR;MIQ4A_&gd]>
Id)0\F+53\6_[/,La/A0>g#eZ^-ORf.S@-[&KC8(2OGKG]6L-S;;^dU@a##KB+GM
:MS6dgX-H(R6SNeKf\-XZ6fK+6g.M78AX<ELGNUK@OZS0\(2@362=BJPQZ.@]CGY
RaY^7(SUH[,2SBU/ABUgC.P5FN]8?F=VYOUSDJZMP(#X3G.dJAO83@;A>]Xg:6C2
/4JWD.1R0A#2H+RC<0MXSgI_@cVJ^gcL]C-VQNQ/0/aYVGR_;R=__@Q\)SeFQ,E;
9+PcAL(3A@=dd2Y25cB6X+gW]&G@eF-N=(M2Y^GgUJda<L:K3ZCSK+3WM,U..+_#
gR3Q:57EYG4\L1YR3B^DTET>UZaLB1727fJ\DLBLES;2BLb>)W31GVOF]\WST8X2
S+dC(XP1SdP2MY](g5^_c-ba4KU,0Qc(<;-.0;Ob766/^8X:-H6L+IYYgC&fRM;]
D5UKGM3G+GHGU<17,ZW;F(&,76R2R06Y)?JRG)Wb76a2PXZ2JYD3WJMSF^#7f1.0
U?=.IF-(4<UHVc;>()Z<WT1UN(:33_C\c,S(\8bgDbJKKTY(8S=4cTY)=,7-6b3e
.V]SM5)>D_dPY5R\Q2(COFHcf9@F2B17)g<4a]f@fb/Rf)S8\)/Naef3\9+^)Yc+
,5FX]5<RCHXc(U^L[KVOE004#2Ee0]H/V/ggRG\[W008H;C_O]cb-V_.c2#DQ7HQ
PNG?5T@5_526-&<_AP1C-(6&AdIOV.8e<IEf9K<=)I]V8H^&>)cW/DZ2M6V/YDJ2
(=Y5KI/fSV^\#TF4][9,-\ITM(=\J&&TJY>?.?dHMH-fdB12a(&9C_Uf^Uf/Fg+7
=K-BNOC#c]DL#Y\.cBK\X:JKKfM].A5(,4\/Y74aX8&c<D-OV7N1J1/f,a]=ESU)
(NQW&OIUO92H_6d[X=NDF\Kd2)O^@T#1<-H6Eg\N.4<99W_V;H2L861CNc3NW1=6
DgDd&BC<D_&);<C])gXM1N.Z31HXH=+O/PD#]TB:#GMWM//b,PAWK[8g\Y[3?>W<
Q)V/>]^&UT-A:N_c4U]9E35<8J\-1@8K1#E^]>U>]<-c9-,#/@[:0A^(#IJOLHH2
E-)NR2UBYBFeaST:NK\+^;=+[.8Ef,(R^B?V,JV\M9?#21&e(BL;XYWbe8Pc6c>X
dD3_TI]_JEcQ3&GXc=FK.2-I:A^OY6,0W4G#15Y>Uc2Xg9K.L#C_J?I[+41B,-Y1
F,.Q66,[;Da=AB:ZM:TS.Kd]R]BI8>D,,44H_)5ED\>(Uae+7[J+BC98P#[F:bZ@
NfRS+ED1@5,B0UZ8F[08^\YV?J0G;cH=#OQHT0F-A1VfR.<OGU=OF>L4TFO7?S<]
3.K^&5+f];c7aIFQ,-5R\&0aO[\9TU/ab)>;?DJB_7^[#6TGd6F<0H0eMT\7R@0?
8@:Pd5XW3W)ZI@]J9aR+H7Z33ZUfD<[f-^<YOV?\-Y9,WfJ/KC]DPEGL?EPRDJ1;
2&L.X>HKf944_7QC//FPeD.AR9.9ABNNb1]5R@4HU,#-^Pd-2U9J39+R@ALVP+.;
c9B?24;XBAKKK.+#38>dFgT:ZH#9(8,;4Z(E#(\28\58[[G]Kd<4:QF7]f&KcfB_
8W6c/HGZL+BB,Z,H[GLa[#Q^)9^3\6#R[3Q.6?2c7,^+@Z-b/[(Md?1Y72[H=UNF
)&B915C]d,FgOY0HC_C9[R4,S94#>9Yb-#Z1:Le=C?7eU@=R.?,)7;49[aDV8&eM
gG7;dM#AUNAf9,=4g<;?[K=?_g4;W_(W8a+ID@,(H_bL:@R9-eMg1(OQW-@eS=J+
X6.>&/B,W6?+QQ)8J2@&6FU,MfIYI?AI3c#2SK5@IQ;N3<@2P8Y6d+T)A\3N>M^@
A_:NV4^.>SI)T=MH.]L/(73DLK-88d.FE5^aY\QfX/Q3DOQ,.KZ\-.Be-(\fS>R&
&(9]_XS,Z.,7/,-C9.2(]0:_4G-F)]/:e.,a/0Y1:a_^<<VRBT6009)I_TY81?;:
9&MJ7GYY,gA&(8gK02b/?;K=J_YW(Q4RACW5c8QKeLPI,aaK#F4)\68Qb4Yb]DS@
:I:-6?7fId7]a]52=b;SMR.<fc;SV0cL,QD&F2?J)0A7/HH_#8daR?f7Z@X@VGS)
IX+XE_PQ,U5V;-R=2b.#R)(+@[N#:-RVbdS/Qg3/HJFUAb-21EeQ_abZc_agfIAM
NHJ]<[G:,^EX>-E8J/FN(L6aHe_b4<PK5[-UYM^NLR-Y6C@Rc3;eIN2g-1(7dI@f
L;7e;<-Td[A-S(283B?8^1LD34XZ+5G]B)&[=(9b8(b+N/=cI]5J=@-/6[3=_8=,
G.P:aS7>HCP=FgTZa-UOb8,OYR-)I,]Pd]4]gW8=\K:3<ZVFbFf,V?+6aT>#\XX3
MU@00e;?@2FOOeVL(07SC?>PeO(-&?:Y4g?+&?b;X>:@g6EK-.86E:9G\(Da9:.&
LHc;P876>RcBH;,e+:7#)O\@A926YMNTKV.L:&4YI84IDIQfg8\G<<Fa@W/Ce(_2
_CJ5G+K\FTO?91S&?CD&3f3E]#-G(E/g8]ENP&g0/,[LU<P2K/#CQd<K6g\9P2BM
@Id.@H&<S#4]JU,\g4:-YOK+P;AZCS3B+d+SK/AN.S#fb=CgY1(bb6AIS7_;2GN1
1fJIAR@,GL_Pc7PLafZe;+971_C7cT?FVa+;NEUAAYXEA]&X/XbQ^aZ39g^Z7#1\
;,K93X8OeXFNOdKV8f&+5VN:G=;&+Te5eVfd?@6OIUU0\bO+7)6#C\QD_+Z:6<\C
-QXeR7;^6[1T1P),2THb#;X(d?(NO0KEWHZ[c8H7Hb)2[\_GF>QC9],8KNgOK90>
Q-]eCQG^V1UOBf(_9#/XZ0Z7C;G?[Q05L3Dc@.J.)9?&3=@UJ-KM&6_5OUJ,7^2&
#QU:FM5)D9+d,f7<U\B5P]KK4K5+]VMS@ZLJ>B]&d,&-T^WY1PX&Zg)OfL8=##=)
_F^8)VI_,+@O\)@O_OKW81L#2OU204;6B\f@71G><CMG4++LE6D6K@d=bg6KaCV6
?3W?E-/(g0[YLGLULC,41<AZ=ZJ-eAI_F+N,4<-#H8<>bCV.P\1(e;Za>\Nd^ZCP
<Z/V=\>53()0&8aNg36\4d=WLZ1f)XW8[=M_4+FB#@0b)f/();60L[#eJV0LJP^O
Y:S(/1:RTY-A<RFIa,\IW13Q+\&N6,PXVe(d<gC#ZgY1=]8.+Rb:5>0;eJ<+1TXL
4&7P2;K#:VCO:3PV#/W[a8a^P#-&2\P=SAF+].UPUAe7W.])aXOB?Q:7:-M^K=#J
OeE4g6TD+&adF&=#8eK^OJ=YY=(PS:/:d/<3\aA)KDU>J1<R=d,N)2g(2D#FBe-&
:^B,-f,dOZR]JP]P=5P:)b&TgVbUd8SI8B0S>174gY0\;G\)?:16]#K=C+7G894;
Yg7Ta\/K]L8S=f.BK#^^LJ//OA^@QIN<X:eVX;.[0Ig8KNegdT#[ZJ>EaK8?)b^C
EZ^;d6;6.A5:d:]?&CO)[<I/G.H9^cgY5@(=K@T(6&^DZ6bIcaY<=H4UVF_TPcZD
9#)0eS=+[0(]5e5b>F^(JM/KMVXbF;USBbRged([KeG2O#5FD;H?6>?9c=@^,V2O
@c9/6EPY\feP(Z9LBI3E-M:3Q+:^?^P?WK\E=6S\Dg+^=Z&-XU4?]4;UU6\:a<Ud
:SW69]\YM?)ZGC/c/=/fMW=SPA>0QB5#B1J0/^\-A+]XTX-Ia=GL625bOGML&Bbf
E[.dDRVdPDLI,S)Kc_b1bZE6a.?Z,2T<;07[XLU+]@gLW[=J?be:J9DJ)E0>DZe2
SQC;/^LcI0aFI]17MbfK,JOd^e1f0bLVF&Q6@SSNH^,R@4Y)=A@[)e<+_^6Qc(O+
?5@3W#+Y:KOB)b0cS3;S-X3SUVgZAFdH,FT7+S.YdM_:O78&::aE[IVJ>OYRG#ZN
]a&R)b./5]e,NfDVM>f+4?\,-W#0BO9Nf)LHc;1B_9c4c\D;-PK?#d2DB=&DMJ__
b@+HJUGJ(Y;OS9L#8e:f837DV_J2FJFM.\:g?>^cL7:WCF([e:Ce;gSg^J8PI5CS
cf6JS0e04?\fgF>F_=)PVZ39P&@U&IY^[)FM?13M9Dd3DB)MEQ8C4.:Q:534R7f7
6,Rg.aMP.e4XA)TCES<f(e2^^>MC,JBIS<\Y0^:E+0(+)ZeOdg5GZ_=QJ)>]VTg(
EMS-F)0\AE07:O0^IJXb^N,I?/8K8;2X\LO8J8A^MK[@D[[6TCIe7>:/:Me-^9V,
_MZZQ=LDOL0Jc8?aP<,1H-:MQATW<\9-=7@@94D/A6YB.CILfU@V/e0R4;1Z])RH
/KF.UL/1B@)@[eMZI9-.N\;(NPKU:_@P-J./g?42MAMP;=^QeQ_,AK]0(T,KUbPG
R@0C^Hc_H29,IEK]Z4\LEDC&8I\S^ALB;=g3PK6EFC#TcUg+RV.+3EFNC4U49WW0
N5Bf-GRgbPU->\KEO]#<AEE-(]eW,KBTgb&)APKEKBND[ND4?AJVI-3,R-#(;WBd
cg#;eICJ<.2O&WTQ(O=MM8<7-8T^_A8XW@+&LV?b>A[dFFB<KB6VOMSKMT[E8F&_
dR+b-R3W,NMg;bLObEV#(9:E9,fK,G.E#T\cdJG\E-f6.\db@]Md@@cF2b[LPLeC
0D=e\b_eQaI259d^bB/M+;)PK,7+=BS&HO>XUea3Z3[J;FDf-VWRfCGK_Q)b1bJR
Z&)J#RJ5QAT(d/RET5a59DU)?g>cB9\\@XZ=4\/]&B>2@0/]&YM+&(AH]T9P,7I1
VWP1CfKcPaNKK4eOY778_QN9Z-K=PJ07cV6WK5F:ACXFM)4,NH;^_MCE?&gaCSG8
,)dTY6A,8cTA:1E<G9^U4+O-A8gHCeP3CfT)&WQ@g?&Wc<163ceSRbX?^38YIgFY
00+LY73JV@P/:);bS>0?TM5Zbc9M:YA0BNG]&+F_gL09,L-/?e/[T8dMSB\I:QN;
a5Ye&0M@Ca0E1.4D\:dV6&&3PAC^#T)^J;LN5_4+N>8(.XY0dZ0EabT4#=8.Ra(9
7G?#d\=,?45??HFgELHLE5b(Z?@eC2EL-F:+:#LRXaI(C_-6/H/:GKb]JTI>THIN
9CZC6&XDNX\1^.M0I54=X/SD/c?R3SWZG2BV.PVMc4FJ^UL[O25MWI<UeC(XL?XF
I@#^C=1Ce&2S4IQU:bWB+e)95KdA9]f\V7M>7AEWAT-H3&_eCM>D/d-c6V;1X01W
(,C>)-8Ab=efULIG0g-+T];:3F087LF+?D9Ugf,\HT90\#<dF=.9?OS^gR4]cJTS
M6LPJDYX.1Z>V7g3Pf504f],@1G:ZL>T[NW19aK]R0@(2W:aaYBX@cBT_94Ge)^1
__LAQ6GDLBMVVX#3b:Y[GXPNWI>P&<97IEQQ+LFc=M>IFC--XPE2Wg@.>eX,QBJ4
K4A)K4cQ.9X(6a)d+I3WV[LY,_IMLDI6MV<:(M;=T)MIE-gLVDB2/1C,9Ua9[DXL
bG4>+B;2X2d>cbG+[=9>QT)+07@EDSBLA^7C[EKIB9LX4/-\KW)&-SU28D-c_E6N
8<S#B(.N^Z.(KfcZY,eE08V[dWYDV(EV?3HBADD?^YP.M3@[a,RfW2NZN/-O;cM0
9ce#M(N+>CS_D99I0Q@\K8C48&Z9CL+W@M?]5?GZf./9gHQ^DNT\FdZBO=db@M&3
#ZLb4&c:@Kc\>bQb70c@X361g@dcUZYL:ZU#g6TV[W@D>GWQCO1Fg.:OF;IS>QEC
[)0C0W/3I3M??6ce2V[2>_JU;V:Xg0NRPU\8+M3-WCQ?H,#7B]Mc#FWVg7A9e?0D
C99W&I?Q[cLL0WV8M@fJ1X#XV@_J53MM2\7aF,f\EYKSXS[^_HQ2UOV^LG7b\:g6
&.a+b@9\b^W?R5I1>+b:#cHGIW9e[a:I26<(O/TR;04\Z=DcRB533-#5N<?[Z7cI
0-@(9#5^Ee<M,K4@.GEYb)a3FPB^00T)MI[70)7X91AMB3XEda)4?8FU7SQ9OLSB
#HgODZXQT4bRN7;8O^V:a,49S6,D&A_?@ZD2M]T/EJ9OX&0geN2#62?0W&(ROHM=
DgUEBZNV\cY-09ND;T.\9a&ADC(7cV5(AAZ=K4Z.OD&,]\e0VZbI2J(c7BQ:L^g2
Ff7UDa#.1T<KQL1fEg6Q7Ha+&b)DDD++V<^b:]_gIKLfCB+;YK0^]JW=X>5OKa]=
?:42dL<X)_R6ER3VfP8]7JI1GJ:Ga[0dJ;4c46UTb8(4,bJ4=OH/3?QSKd0?^eE0
&VJd;bKV;_K43a_(aHaV9_fRAWU)-#SUC=HN+J03H9N2(>#B;OHH04#[4>H&S(eQ
U6YK&_B/;RY2S_.PI/?A>:g_AMSV2CJS<PfR4RR+4.Qg2]9X?6SOAM-;-/A>fCH2
(ObP\5Ne,0C1[^+W=4OCEOY:AKaO]aW/HY#2bZ8>+V)B\BIA^N:#HHG/NLJ-._UQ
^^7TI1cQ4f#C_KM7F<eL&\F/Q5AO->2V3(];Y(#7dY)(1,U[_&?>G1Dcg4-PL@OO
94;;16^&FH/F+H)ce-(A5O<^3bL/X:^>e+d:&RJa;-D;OQdNESfZY;X)G,N5\]b4
3\T8=PA,Y=VUOP(W2<G\GFB:?GbU/3_gX1I1PG[Nc<N?+c3DgJSD>K^0OQ8bD^?V
#@0fb]T0K4]LCM2b?7gb-GCEU/,;(ZZN\W[5L:U.@4Xc+dD(]MX=1=(Z=d?M)B3Q
?NJI;CFM^;g#=HVeb4J7@4dWJePMOEMA&K3EVZPPUcT6@UaUMb15]6X.Z=6e\:fX
24>[f(;aNY@,]@231#VC?6\1L19BVF@F>9/C@G<J[8LUbBfA1K<MTL?d@g5[W=2P
S/:GI05a+(<FN1QL[\=_VV-e_>=eDbSBHgPd_O7Gc6D9:JU<JgD.C_@XBN9@-U3d
64J2J7861Q[L2fS1][:>ZcR4L4_agHIg7HT+4=8<2g@62K=/?^<^MOaKG#\Fa+=8
#Ea4GU-Q(GSRGQa#>d97DEcL&7Y6J2V>WG)8-FaW&3S8)NQT;Z+@,G.=7,519-//
5EOeD4#eRXV[BO;BZUH[S[QaM5>A([+F9ed8T2E0V)9[>X\2NIf6Z=(F+?8@@DM>
GL5ZO:<D.^)>/?U:28d56bfYB9,CQ,[=4SDNY3=#b4@R(;ON5E^NOGS\b)#(fR<-
I3?EU1B[O^\DI0H9?R&Q#Rf_W1ZPA7Kd1#A,L5XU1PBHNd#fWBP8g8Vf>\Tc0:V9
U?aEb3[@1R\?EF^eJe5Gfb4eI<;.7=S2?I7-=@V)C2(49AY#+]);VKQXcOX7WF(Y
ZbY,:Q#R=M^E:@EY0eO+eVD+8>eV>RBK=W1;A;:_A.Rcf4@.eNM/g)J[)XO0Qg5:
)f^<:cQM/0ZH(fIC;])C:M@D)XNH)S@MBe^Td-U-gK9W,+K9A^(/4Ud>\40O>_b)
g8T#fG78Z[eN@5d5=#-Fg9>cW\a>_@fO,KbG9,&Q=fBE6FIOVCe>\O/d]^fWR^FS
e.ZE8e=6_>_WW+1HCI<c[WTT9Y)]NMQGg:&ZQ.\=B#Of/Mcb5OK2BYDCJ;AH4&F-
)PNbTST+ARb>c9#ER@af(YR&J4Sf#8b:CT.\Zb8B2J>.73MLXCD4d6+H(LI3-37P
#&P0)V1_\<X,5(=:,P[V;]_383Z-J@)BT[>_5HC;,)T/W098X,<g:ZdZ2<WK]5UW
C:V@^H3J)TV\&^-fdP4Pc86;&Jb=D0_Q=]fg3-#+FUE;5J;875AgVO\G6;.G4<DE
^eOfL&3[(bKI\S\BEEM[O;Q\=J?7NFK\7S+#[]7LZcX?TFSea0U[6dCLIGb]&@bd
)Cd22Z@1Z?VGdRS.DWP(54+7288+8f(3fXCSPfVAIC0Q>gOM7FQHZWAN9((&V3-D
Q@&31&<6NY0YfQ#LM:[:@6CE0/>FW7>&FR7eN0#WRO2fO9&.2IEXT;KJ@8761JWQ
38^#c6O_+E+D&d]S_41IBCP+2#DS.6B5=3;K]<SWXaMGE&Y]P2;-=SL-HHXT>J?S
d;d[_-CZTTG<X9)040e#>FD^^N+:g>@gL=,b1MEGWIHX+=[+.c<&QI9Be8E+XUDb
^?g5EbQ_^WT+XTPA\H?@X):>ca-SJ^Jb7S):WG&V,e#OMfcdGDUD]26Ec?2V1-P/
)\aZLW)5?D6()<L5NH#<0BQA\<.VaT6<9UQ4</gdL9\J=)?g@b@=PH/Ie479/V9]
IbZVZ>c>:4&TdAOJ83YZDE[Bc;:,>6_ZL9)Sa>gB1-4Ya/AOPeb3HH?gJ(L<9Q(J
b[]GQ33F5SX200JF3]CZB]?M-;[CI+bIMU&T9dB@8,Q^KZ)E/S,2L#X[XJ.gPZ#?
N(D0Kfg1T]ZZG6d,.VGV#&U.N+^c+b^#F171TW=V90&BK+e:aRc+f,#Yda.K[_W)
d/X1f.g,[eZM1I->Ua+2^,-2Bf0;<2bS\GF9VW@(QSY3=1NSdRFDVWK\KZGg2,QN
T[;LKH[,,AAAD_M]8=Q2[191_9/+OT+>5UBH>gL>?e1-2VHcV^Q;#UFf[ZeB+RKG
DG5316(DfeF9G+-1[g>M:=7d[<0A4,H)2Ve^+)ZLN;&ScGMc&4c]+W6f9I@64>;B
X<4_5JHa);)MG5ZQB:H^IdSc).K@[=SN\9YeUWH^d4A<J\?ID?aDL\aP<Ra;[?)@
eA3S:YRCUB9+c_C7Tfd0MgIPYS\?/f;3TNS9QMae[6D1U814A)bQJ-.cNc^P8@@5
fTS#MR3UXQY@73]<@RQ?\SH0ba)+O.&Qf=11=[dUSY)S:YGO-9+bS7V;9.3eL4KP
5VGD#PHX;e[Sac)]W:H-ECbG6fcW;GAJIVF4P1@?-0a^3ADQ59U?U7<JeF,&d4IB
2C<\Z7?g24VS>__2\6[OFMLQ7[Td,,SGH@,Pd(fL^0/V^Cca7YWJ8(P9-7XOaR#7
O8a7M1-8G,-cEaK390DGAM=a=_3\:8eTF25b3+b]V_e]TKJBc>8cM7OQM@T/B9-f
TK(fO:KgCU1GR)-3d#@;KS)PIGWcV@VDd?-c3#(-bT;)#NE6NF3HFHXfYe5fBVB9
-SZ/fae;,_,L_=RWc4E6-B_KKR,DGLMaP>K6fM-NEd?4?7_#-AQIg-X?Rf9_>\X@
8b6\.\be9#\\Ee[[[;C:c0(L+6MGH>(f,=L9JMI:P<Q,](U/Jf^g_:9SUL/PbBf>
K.YS_a2]>^BU\aT)G7[@Xc.S_EUYa+\W3I^<QDB;Ab@)69M:.<9;X-,EaYb86c0d
4\VVcdNS[g5?;POQL-M]+SG2N_DY=Q9+Kg-5&G^d8U.E_a>7aI0I@=Q6A8JVR0R3
cPE3>&2cTR/[(ZLQN(,V5I:5-9F[\a/I(L8fM;D3G7L^^OW(TA4=K#R9\XbUW84D
K;V&>7&;WG<Ib-?;dS\GX;K(]Ze-WfE.9TLJ==H7CAc?Y(]f<cXZ.?XQP=ER7/bf
J0a9f>_F4g;6;OADSR\E^6#BYN<R1.+4]PgF<>eO98bX<[_ZLd<N8J>;-YdQ2e?b
&9WC?)WR.&D]+W=O5Q_:)P5?c0[&O^-;XKa]5]:17(b.M_24C\XIPA^,&U/JO7J^
LKOGca)Dg#EA9BP+cFOLPg\E_@K0CH/JBL4+[aK[PKW=7eK9(=c?>>Xg-1[Z:LTL
\TQfSN>#7Bc+:W8eX:90.=4?#+,(WJS(;e&A/aD0MSf4JbF4YT3a?\3UX4f[KZ0J
Ca_a/#;=>^2)@R]:[I1ZR&:3FH?Q7=9&N62[:7RSL?X]_d\0?(cbF<8TOI#NPU];
.9GM,#^NOYWeCAYHME<()e,&_^X?A>0]2[REK3:ZK2<.@B(,4.SW-H3HHT5@e5-A
X0FV#OJ;?0XAL1??8@2aC_&,4[31_OSe^T2:/XV^,GMc6ZcKX=(Z6X?H)\QS=3a[
&[B;Ub/I45_5)Pc4_D(NY_Ja5D0V2O5L-TTY@O(@cE:RD^N03:^cAZ])#d5G\=;>
9+G3H^cVM5B)\4#LaW-,d?=0UEb=;_Hff=#Uf>AT0E0<QSab0I&?dR;EJV__Z_F0
;@_<_8O]EDNB7b=EB-_@I8>=+3\YB+X)&IHN25PE8O->>(VWXW83V7(]A\.[RW++
XBG?eP,-@S(UY-Y.WcPCdUL0(@A2f)IVH@M(Ia==&eC=&c-N]UQdJa--T[P)FaHK
[:]7.U@/GWc97L-eb(38b#IC:^SR8]P=L,[B5;(#(7S5bcMX<8]g-d<HG]H@2\=&
eJ8cbA_N_6Ef/4aV]9:8aG5][(dOOQ-ANQ)L(S-NSB.,)6AN)c?/-TCH:>TPPSQ@
f^GD&3Y)[O&>RK?FfcGaacL\-4cQ9[?cXcFbN,NcKT1JUKdIK4854NcBgcW_;C=>
@Ue3\.RM6##+?LgPZ=?@/;d7)FHfLF+c+f)B1N[H5S7@(6OPI)O?S+BL#I-@/I+a
R36(#-E^WKZ5MgI\MEL2,?E[ZAP0YQN2LDS+^)K:0L=N11PS:&df__>LLT+g^Q;3
;N>LgV&?M&W]QXf9UIB:a.&C\J8,T3^,B.7dKYYX>NDU)Z/BCK>&7-9.@8Ya&d(<
4Af1^e_GG.H+3\EU#c@>(McB452]I0KN4VNK2W8@V2@3PI:d1/R>)Caeg)34E=GT
;Uf[4eD@a@,VacFSD3R_RT6aR,IC^^FQaE_Z(/=\f&PA=#b9aDSS^0:F@IaSg@_9
Y?S9=#8NY5)O0H5fO41&J<Q[/72IBLVD10YbJKLcCWRJ]a=e/8V8)=3e^#+W6LUe
J-CD>1;FT[0e=<ZI>/U=7ZMW(I8KQW&3UN/e]D4J9QB6+Z_-().1:IT9dQcR=9Bd
C2K#L?5S_@_bD.(?KZBa@9=9(e\Z(@H.ON<bC;(X3^/FD3=2f1Se5ZN_DN^8UaOQ
)FDV#QVJCKSTY04SFF6TQ9>@b4eBE8-G<E:Q5#S?P=/LQL:E@Ygf@=JDR3&BIIC\
C8>J]9GGY;9W.=G.fgZ7;<I70f;8ZWBJH)9Q()(+]=NVgG.6K<]X]CB^+-VN\NJ8
T8)aRV)94e<&dYgP)JZ3>+OE)S4^AZG4Sf[S/ACOe,/KGbPYIb0BC7H.Zc#99R\@
b1\<<(AZVca^SXa=a&0IBc;S<d&SE)P4+(?Tf1&Y:SQUfcHa\a.9YL[9YUIZS61]
&AAWdSC,PZULMcgDK/>>Z#7fNe&MT:,,_6P^;7+(aI;@2GEZR2=d.[Q?3#g,?8)I
cfV6_5KOH[3F9[C0/X6_Z[R:/=(>7T:J()4OIG()C(<1gY:[^_6GVb>-=FATVada
X9VB.1VHS&]C?ZGb347=I6&?^eU&19>FSYE?1-K.Af\>@5?==2B8)(;&[d&6V=>7
XXcK\:-<0\A+Y\cd.@d0HA(XZba7eb1Q<d0_8df#43cSE\SRI0+(;b__@T;G(BgH
bTDF>JJ0D8+,_&)^._BU90N6[8O<QGRS.N3E<W_&^T.S&f]EedNRE_fA>bB7Wc:D
gc[H?X#-D5GC@8R^0C(DB.BgRP]@cA?^fG=6D=eKR@-,)dI.VEJ>/UJdD0K2SP\>
2U[VOWf(E7CQ:D\(RJ70Y(9MfUH5Y19e.\11,A/#d5#F8ZH2):GJd>#gd7HJUF_6
:5ed[@CJF:e\J:FP8&W47YM?[(]]TMebbHPL4W4:bRRY2^dKV60LJT@C;<[/-eD9
D^LOC-G73[b+Yc;(;=65/QGK&.:(b4a^?1958)PBPB^]QeG6fMSN[X=2;G-(2_1:
+_F6a?JF(W)_+:>>&U6eIOOYNML?Z/AXa&0:-N1AH(F>^a)b5/aE#T2]CS?;-6K?
[-ca^^S(Bd)ACW;LYZ<c^S1JbCb)PDB4QHGa8ASHYM/SCRNHBZH?PBf9d,J=JEF7
#61LQ+/:d<3#K;(VZ32O3>^QFR:&F@Og3:aH<.[dMf8+#e4AV=cF3J2OaKH54b8-
^&NZO&U?g1[7@QCdTb^U<Eg<_1(N_<+/gNd+6f&T3c7(7cL)W7?gRc=4C4cICU81
PNcZ;9)cb0FBeAg91[9HE+HOf.D]:97]^@&R6HJc4>Z+0F+\PF\,dAI,F_A_gFVg
HJ)ZN)E)3L^6[;P.HGJ7.Z5]ZSed>S01KOQUNL91O,FAH4UbQ:Pc^W;?^ZV)D7I@
@D/Q7.0=N<NXE4S9F[]N-+aC_G=:3AMPKQM9He9M7FVQU3dCb=>;UV_AA65ZNf&&
+?Y)^-V7.&BK8>fPT3V;#+P@=\&\MgP[F(a1SOE<IPS:e)>CVZcC^2Z)Q@@N88]2
U#^eg?/?W7F3_4^C)-G4e:XO^E[/M;EUBIbLaWf]:4(UDaa?MK_fEJ?1c1-:;7O@
/)]Q)C:QT]Cb6(fFKYJ,d(dMaW/;>+<b&ARI@2BLbH;f:>d;::TR\Z4Y)YM-Y0X.
6U&ENB&2K?F=+d>@ZH)]^DL@/If)I>e_GMEISO1&\GAV^IW(1+9>\4>gX77cfGA/
AG7-3ZCZLaT,@VYb@BDMUVY_Y/LPJ5?7^=_/K4C>X54&NW0,Z#E\JNaQ9M1\We3U
fe[HB:eO_D#g95A4>?2@Df5J[Y6#/-EDZ<\L\A0]9fS^7K<Eg,4gF<;+f(#dJ2+?
WY45L<\)GA_B2ODT[BV8T;e8_:&Ne4ObOQE.ML,E=4/]7N<&c.&6YUJgSfU4)7^(
,UZ-_B5O8_#0N>[[IHCZ2:D(;]30GUD8C@8M]K7-ZX/c&KSC;I8(E7?1RMWDQB]W
^[:e@P>.eBH[W:^:]F+)3F(Y3&3/9I6)D\+WLD,3@f<#^E^=L]_7YZSSLPCRPQZ.
b16+\G(OAe.aUdd;,DA^OLTgU;N83bL<e1S8HMHT]65c(\N5ReJN(44#[D?0.@KH
S;^TF6=@8;@US=#F0-Z7W/0>W74_.KM:?H3@T7fg3<IKdM8/T#5G8@3D0PBTCBUD
g&309O9D#BAUWbeA(O<FWP@S=e+,&K3;2GIOM3E9D\]_H(CH/_I,S;+J9_C)-Z<d
@R4eObgR;/OM(HSg.M2.&&8,d35e(A>(N^)26MDX0AD3^=+Z&E674FZ-6I6_YITa
HGgBW./41@f,9KF]_XPP:_Z.^cI9Z]G[>8)FbZg0/eg4L6d7#7R@P[N49V_3^P5\
08::JP@bT?-POS7TVL:5W;BS^^(5bXJCFH=9?_/c\cU]HPOgd,^6=UY?+BTT3fAP
JL^1A<TTJ+6g2,EBP69?O^fP^BQOT;D(113F&d_bY[GeIGH.QL#g>G8Cef.6c@8D
QCV;4RK)3&MCG76?J#Y<\&(AMg,7J&Z7Q2aISS?]MXX&2O;;O._421MI0TV^NZ2e
\-P1b1;Q2JRFK0\+>+HaXB-)BgELXR:]?W124@1VUKVW8Qb7aN/e]U/RXf>8Zg;H
+[5]V^-,53V9fV4;[F(BXE)E7H3,g491W\PV-bG5aLA);HLI8P^U/MegCMcX#/c+
<IHZ>I:XYc)(U)88NE76TWVf)aU#>cKPUS9d[:<64[E)-KW-&F84J2)8(gTQ\I^0
:2:84.E(OWVW)3cTfH\WOYTX7Wa^fO]+U,A?QQ+U+Vg<8ET+Ie>>T_WH@eZA;L-;
P7]_]536QaBI1GNAH81AJTQ]9/bUV,7aGC08WX=.#a<U:J<W#SbV?3aGRJ:CJDI/
:]LFe9LJKF#OU(^=#>V6\,<&cefQ^5e815fA+.@0[KEd/W9K2bY8&Y)TZfgg(UG8
E]>C6JCHKb);5/3/_>#9XDL>,7KBLBW#2aN3^#Jf#?S;fD\P_]AZK7FS0K#2ac6f
bM)>;EDD.Ag]8=3J6&f?W7#L?B>QKP<B3a81K7,]T2@GF:,X^acY-UJV>]FEAGaS
FdE0P-^_;ES=<4WfB-58_F0\AdJd)[/50_;dIb53,UF95PTPW<\:P\P76@MMfHcc
H;C_U+KF2f&5.=V_]-507eDP5B3=&&ZgKY(gC].g7E9Z5W5L7?D1;NU7J61?8ALT
_Y0B_CK1U</;QFTI=;S=Y];cbUH@]aX@U68XfO0]SMZ1&a3-UZ^7(0a:<^HfI]..
+Y[Jc6-0>QPG+_JTffB=,4,^2-W.]+Ze]M<9S<e.&X&cJ,X].@V(IAVXGAOUP&[_
Y\3Z23C)3L#6TL.7[6/&P]AR08,SU?Z)W-@c?TJ/5^5cgU9_K,;.U?XbRK6#=/RX
FI+R:8,6W@TR9@^5(SDA\>H_eUC-G[([4A,AM(HEMT2J+X/f.UM3ZK4KgVYKPQ^R
ABT[f7\D>(2F-E-cZ7\CQECS]BMB35ZGaUZ&W#996c3:ND-NH38+=@K+>]f,)KN>
12;VM;27+E@f[SW4dA+IJObXK7=Q&8Y4,Q9W<8?bY9Sg5\&#1<HAZH[T99]3SL&P
CF1\GGV/)DZ([e\+:1E/<L];Z1=HL#0@fd4769DJQY67K<P7WT=WF<b&]?@W<)(2
13:-RVOf=&6fR@(ZT&#.H9QIS#US]e5DEINXO8>ddJ9S[e9f#-+7d;f&Wb/V[D2[
A_&7.2IBYAZWHAdMeXW]8c_T1QE9//U<Y,KX_UN?J+=P8M4g[5W:-7+T]+928(;=
RM:,Lb>D\OX^Tc9\AY6)QE2gc3a@\&(JNNHd=\[b.BLb.OgVS,VN)(ZBaLQ:V(KP
#cH-#8+3#L:P,O&2#8N.CgU;F:aZH<F0@^NIJ3SL]4agM.-ZMDeT2KOf^+?g.P9Z
(f&P&7GV8E3[-7Z@5DW6c+FB4[--[\5.O)YgIHW28[\bH\+e+]a,UGJ]/?XM=X^,
#.CY:6UJ;X&(9A_IX)H;1JccQO5BfV6BaWO2C8ECN-_J8#aW/8UP]bMI[52<AY23
H_YZRP39fGgC,FM8aNYH_S15K>[/Pa3633L&J141gYYd@R<=e4+.N)6c=DB9ZZKF
[c8aMg,?.4.4U678(eOI;\e0bK=+11EF)I-ee@a4UXE8aQ&8cN],9d4G)V\&1cXU
Y<Ca4/A=<cQS;Q59LeLC45-N86MJRN74eFHX(TF56Y[YF5IS):UX/W4\ZHe?f0&M
C6&DDFGT<V_b;36P5ARW\-)gVF.8243K,AAX3T]V;F20C:@:RO0fPV@PQ\J2@]1U
V/=&-3]Y=0]X]YaOS0=R37Z4DS.S#84H8ZFB]N3a.EH&RC>+#E@:gZ-\<dK\E<&\
TL.),4b6eU&S(7A&JY@6MdBY^N4=&H^dC8b_UUDPT=gPf+SH@-2ZD61T;)V[G7a;
<A0<U;Y#8O;+RAa=1Kd\(]1@=#.c]UGFI2@</4BU6g.<?XL4]:KUVI^Sc9\KHD:F
1E11aHWHD,RN)96,A8b?QR<bO,HN/:adZ0eSQIc)W/MW(U<^]4NfN4&fW=RG;HXP
EG)A5+g[Bg=D=_O=e#KcEY_PLW?/<Y=VW#e3@D6#aU&GNC52CdLX&1WWGf\(b<eX
AP3X4SE.O9#:,;K#c9N>+K,IO6:<^fWVRJ5TC(13<?I_8CXL::?2+45@W07#P0;Q
aE#2>7]8#fDPC+33gYMMK9,I7$
`endprotected

