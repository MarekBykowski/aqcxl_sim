`protected
L-@[EN^J2KJ:]GQcSCgM/[Re1AEXR^Re,2BW5C@<=_2X@J->+NeR1)^8Vc97KI,#
-+EE+5@VG\[[_S=eC,NX&8L6-=0JROYB]c?1(VE-#PcC11RZScP-G>:^RX[]RDgE
dc.O_-Mc^>gX+McX->b4#06V5JDS7(TAGE?a,0D[\KYNO/9^.K.[?X:.)>A2-FJK
W6.+bdJKQ1Rc=D7Ig6VI9OeZ>NXO;];Q@$
`endprotected
`include "qemu_enum.svh"
`protected
?S8(<Y.Q0G;Agb^X^5VJ4IYbPcH9WJH/@ZD@2&dCGaI8OJ24Y;&N3)SC_=a0@#Ba
,b:&L+:^XUG0]-[V,afX/eM+W:dY:T&2YVJ308>&ZFAN)0\YK^6g^6]\U9e<0N.0
-fP#IN9=aD3-3gM;TGTB-)1SGP(f&L6/BJ&(P?X/PLV&JTFLW#)@1FBW.62Y,0Z>
c;(V5W_Md[F@b,?2X/NE=M;FW:6g-1KDWeMVXg@4V6-Rbc77V/@IJL<2TR818YV<
CO-\06b39.M5XR9<35G:dT7Qe89,/.Q^\6,/K^[3^EKSdPJ<8#J0gTeH<A(gJPC8
gQ4A78X)Y7S\UaC6E@fNQ@^4VMaHdDg+c04\ZX[EY4&[LJ6NL:8[M0M08b&H_1]_
KNM9a]5@S3-]5c0N\,DBHgT+CCB_>)D@JbAGD6;f1?9\NU[?9E<G<PHG=)&J,AY9
BGc_Fe.gJUIA66Y1R,K;QA,&6d[/DK6AJYX-37g??/)55LbP4;Ddf6eYLSVD_GA-
E@TZ\Z49\RN71D^[P<?EZccN@##T..g_9U0,IWb:7;=I8Egf:Qa7Z.WY9gW^4#M4
d:(\CNRYdC[^+F(VAH45?G\6Sc9>e<Y)dD9cN96(&Z/f9AE4gAcJL_>YFS0B>g#B
>7C\B<\ECNAGY70(faB<G2=YV<ED^AVM#0+-)SJP)I7HWAU>O3G[8^U]Q)09^[g]R$
`endprotected

