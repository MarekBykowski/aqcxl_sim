package qemu_rx_pkg;
import avery_pkg::*;
import apci_pkg::*;
import apci_pkg_test::*;
import qemu_simc_pkg::*;

`include "qemu_enum.svh"
`ifdef INTEL_IOSF
`include "qemu_iosf.svh"
`endif
`ifdef AVERY_SPDM
`include "spdm_dpi.svh"
`endif

bit RST_TYPE = 0; // 1 for Hot 0 for Warm/Cold reset
bit PM_SUP = 0; // 1 for Power Management support
typedef bit[31:0] payload_t[$];
typedef apci_tlp acpi_tlp_q_t[$];
typedef payload_t addr_payload_hash_t[bit [63:0]];
typedef acpi_tlp_q_t addr_dropped_cpld_hash_t[bit [63:0]];
// size in bytes of the simcluster buffer
bit [31:0] qemu_debug_g= 3;
bit [31:0] vip_type_g= 0;
bit edb_logerror_jump_g= 0;
apci_tlp dropped_cpld_q[$];
addr_dropped_cpld_hash_t mrd_dropped_cpld_tlp;
addr_payload_hash_t mrd_dropped_cpld_payload;
bit[63 :0]  _all_one_64 = '1;
bit[63 :0]  _all_zero_64 = '0;
apci_atc_mgr atc_mgr;
bit[63:0] ats_xaddr;
bit[127:0] base_limit_Q[$];
bit[3:0] evict_mode = 4'b0011;
bit[63:0] max_clines = 8;
bit[11:0] pm_cap;
bit[11:0] exp_cap;
// Do not refactor PERST_N this is for sideband
bit PERST_N = 1; // active low
apci_device ep0;
apci_device all_bfms[$];
// use integer instead of int to avoid vpi issue
static integer aqemu_int1, aqemu_int3;

string sc_key= append_key_after_user(`simcluster_QEMU_key);
string edb_key= append_key_after_user(`simcluster_EDB_key);
`define SUBCMD_SHIFT (8)
`define CMD_MASK (8'hf)

`ifndef APCI_MPORT
`define PORT_NUM 1
`else
`define PORT_NUM 2
`endif

task automatic set_hdm_range(ref apci_device bfm);
    apci_bdf_t        hdm_bdf[`PORT_NUM];
    apci_addr_range_t hdm_ranges[`PORT_NUM][$];
    bit[63:0] ig = (1 << (8 + 6)); // 6 : 16 KB
    bit[63:0] iw = `PORT_NUM;
    bit[63:0] hdm_base = 64'h1_9000_0000;
    bit[63:0] hdm_len = 64'h0_4000_0000;

`ifdef AVERY_CXL_1_1
    hdm_bdf[0]  = 'h000;
`else
    for (int i = 0; i < `PORT_NUM; i++)
        hdm_bdf[i]  = (i + 1) * 'h100;
`endif

    /* Create RC HDM bkdoor mapping for single, 
     1 decoder 2 ep +APCI_MPORT
     2 decoder 2 ep +APCI_MPORT +SEPARATE_EP */
    if (`PORT_NUM == 1) begin
        apci_addr_range_t range;
        range.base = 64'h1_9000_0000;
        range.len =  64'h2000_0000;
        hdm_ranges[0].push_back(range);
    	bfm.cxl_bkdoor_add_hdm(0, hdm_ranges[0], hdm_bdf[0]);
    end
`ifdef SEPARATE_EP
    // for separate devices
    for (longint i = 0; i < `PORT_NUM; i++) begin
        apci_addr_range_t range;
        range.base = 64'h1_9000_0000 + 'h2000_0000 * i;
        range.len =  64'h2000_0000;
        hdm_ranges[i].push_back(range);
    end

    for (longint i = 0; i < `PORT_NUM; i++) begin
    	bfm.cxl_bkdoor_add_hdm(i, hdm_ranges[i], hdm_bdf[i]);
    end
`else
`ifdef APCI_MPORT
    // For iw == 2
    for (longint i = 0; i < (hdm_len / ig); i++) begin
        apci_addr_range_t range;
        range.base = hdm_base + i * ig;
        range.len = ig;
        hdm_ranges[(i % iw)].push_back(range);
    end
    for (int i = 0; i < `PORT_NUM; i++)
        bfm.cxl_bkdoor_add_hdm(i % iw, hdm_ranges[(i % iw)], hdm_bdf[(i % iw)]);
`endif // APCI_MPORT
`endif // SEPARATE_EP
endtask

`protect
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_2)
//pragma protect key_method=RSA
//pragma protect key_block
AFUWe+h6bJH4dGToJYy61JDIfdAbVPBI26f9dsJxBCsH5c9YJtAAlNTs9FpREeRW
Q4Oxkiv7nLvdn4Lr/+mVZIXPFeliT6ZofrMgB+77sgEl2ts8tksEscz8wXAU8R7l
wzKJx4XMRw1ZcAcfXxJRrCxs6TLlOX0+o4u+c8l4ojnBhVZuBBJWXQN5HQP0qxS/
9Wx6QrTDxP9nIEnSmCRjT+3R+Ov4NcJt17/aeu42Mit7+HzRwtZXGcUqjZ9apVKw
MSDp7fwiLtx/r8vTpnIO1sgyCvd/HKYb96teWXKdGTusBtvJdecNvsagsYS8nhj/
syVFDkrQ8H6pF6XlPWs+nw==
//pragma protect end_key_block
//pragma protect digest_block
pGLWamJoyk87FZ0YnmcqWjQFUhU=
//pragma protect end_digest_block
//pragma protect data_block
1Qd1B8ZEHkjuuBh6YeTNjEkLN66ZbN7cRQM+OuPPCAJQNWXkrTkJzLZnn6GakT4e
f23IypCprd+GCZMXwxKIdFGxeMZ7PKFNCBew3QXiRRkRL66RuSPncb6FxpI+tN5F
5galiAA3PRuDTIl+n6FdtFDroGr/IEuTzOZeuSTi4u4eG4aDai4XQsYzuYmapPl2
a/pQzSOqtu4Oht0At4f+nT9lbkO8jnntRizW2fzxa/VVJ0T9TpQyJxyuNbTGAvjs
XTiYyybGy1zmHAX9XBGCZoQmOQ1iraVYGkhMRqDcW+UuxaA48hMz/CloqOedexfM
tHCO+fiFgJCptLh10prE5Vc5FTkSRlBlunQHtGNfJ2tj1CnJ1i0MjYach2WsXgMV
o5F54H2UTgFuh8jIAKUean2aLRfffOIGH3w7C+z+Oi/4rgQ1fwRqbR0wgjPvmOxA
DCRe0tA9ZFO4SyRPs1xBYytqWUzNkHDVFdiKkhY6dFKj8T9ZvaGp0jeYUh2i6n38
m8e9NBXoP51FbvsBcWdKYxqE0gyTXI2/MmB3+KQv+55/rUaegUKqt5xhbTpjz8A5
U6TdqV8RwRAqB0WZz0ATiykQwyNiUETaXaCpAO6AKQSZHSFyhOl89zXgSb+jvYJ0
UKuaV2oQyouyvtUE8gAGX50Qfc9WemyvcbuyD+v17W39eUpGenjX52DKa4+qaMzl
EYVFsqQVtvZBf5LY+RW2rHLubxrXYAcCmOPcJZl7zS8sO/q5kIDdooMl5fXgV4Or
O/DlagoFhioKsHyf2m+2VM0e1yP9oYnHuBQhukByTlwKMpXIGZQXI4r1rftSFxjj
jJ3SWg70DUdXuzfcMC3dIvqPNzgrfk57JyFNTpPVAoZ2hOGZVziPyjPSP34FwbuC
BammrGAoIKnytAfWF0pD6T6XMvexColFPJnwawTYExiMQa85hy4zTI4pXzahSyLq
mZ6TVLLi/wbdW+CE9ChzJdhUh1HNVYz7Gwi63BNucb0TgfkCnEqC8V0gpW/viZ08
KhWI/ebKIxhiS1lLJZi7pcf2+v7FBU2M6xySL1DXbxdLJsekj/d3k+sSNuTg74+j
n/7WNMci7qU8Isg2XmZzwj3KM/kDD+ehN9XqN5lpF7FKnp9lys6PutK8LwdrE1p4
4us/KTzg/JxX2gZe3cJz7ENR1fk8uP4RGmeYSZIp8CLcpyh0vKrhoBOBgAmbg4Ls
0aaDGnhjG/EzUDvPlg8fZ1JKlGrfPrOFqxSnLqP64wFKUB7HcrGdq+iLJEZy9VXi
RkRhGBOz56Cyp3QKyQBMutZQuUdbVLAA/JY7BIhHjUn2W/q2MLjFrV9iE3s7EG0/
xD/iBqn3NckbD/OxPp+Kk7q7lZu5TEuLtDxLf9tCvqDNo/6ibLAuER5i5aK2B39h
ZaHxEbXrsKbPz1+Cly1B07vXJ8q1Z2LCh+cxigkWukUkP/c2eMhLl/jKI+Czb2xv
VWD90FtwRiXmZSRDASiGFCsQW0vXn/fE8jv6687x4fUvNjEiZ9udFg/0UqSaT9T9
F8PLHHH1na046uxsB9oGVcue3WDpGmuUV63TGm5e57gJcStN9yVmyK3fXyGcq2Si
HsYXg4cIMnoJOzu/J8ie+ilX1cd/THtI2JTMLxKUWtpKI/M4JN4Fv3NvTmC+E+ke
0PzItp9uCpQ/sOLwgRz5UuuP6s0zgfhCyCpCtj0ev0kJDVI59QN9UhlclxGjIGIU
KthgwJ/Jsh7DgREU5UKYmRS4dpO4/cZr0pMvjfLXVYvoAGpBNksmBHdxCCbb7ER1
TsmuySX9w4VPDhEPkCGdcMUx1tXmsbdJdMGndYtpu2lH2EsurfjxlNl1WIqX0EFW
TvJBU/dsYC8jf9chqoSqOJAe3FRo3aS+cgb3p8QmZqzvfmAweEFXU7WdGh0X92hG
a5y7141cfP1rLm9rZ3/L/vVkN2/Bk6WDXxEvNkaiubKWAC40R4Nf0wmRuIW3MXXr
4IxSaYzAQDNz1+N2MP/t3WZMyLpb6QBkUzoVdLeagxXiRtu+k48rDEosJJdZVoWB
s8SBvBDT/9akZv4qXUG2+SJYQH32O758yS0eT2vnookBDE+kaqIFaBaP1DluHDam
EC5qveUHTI3K3m6lddtBvNWSS9vtmnxm7g7s2X25xCQuLsZI13qgJxiHqqMlxrwt
c8487J4wnSMqFOW1EuUfe3O6i6NNOdvHCc2ZQBbkIUrqxTfgwSx5EqsZCbDl47GH
uaDmWuH5xHBq+FEe78OH4nRGmYsybEhlYgY4Z7x5d6GVq83sEgisdHIJnSgtZXeR
QryISkQw2xfwhY6yP7d0MxbcJ0/EnuYkGVDBxXSCxy4wxYBnqn/fdpi/cVCFUQtI
aNutbdOwqiEt6MM0XXgeMRxxOsRQMq68Ic3RhjKbULCMc9ELecpDA1qhbyPfWSY+
hpkfnNceYU87LlqmrdULsKCNmZkzEgE4SatI738aefrqs6ZZxhVX1GrO3Kq1rmv3
fm5p3KTaONwCvNzXJQFuXQYXf+9D6RFeRXeVseb85jtCx9OHef8M2DSM/uIMdGT/
TH38cWMZO3uzo6SyRMhsoA5f/Q6z/k24SBeYPkw2gV3ampBpsFp+E3SAY/RjBeEq
HZ1ovEtys8Vu1ZiC9w5d3lPWpgYQsO2MKXapQOBjjJe8txlpmyQ8iK5Lv7QKDd28
upvwBY6VBvA3iuATLQMWsF04CuSn7ahtAv0crLqnGlzBqELDvOw6iR/gpIbH3qQ2
2QjhprqOFgBX/a3EXO3XKh2sE+PQ2k0rJ1bqahE7sy2CaG9hUrvSAgqhBDu7OmYi
CqvyuJlUkxr9Fvqqbd1GszoidUPh1kB01f8/aekrpOQgvP3HUe0bJl8z0JRwo7hA
DDFkfLe6J5laSAamGVZdCpQL7tdccLbnEh3eruRSQEIsVMUb/b0S2cZmiLDu81p2
i1n7H+fAKKMOuVULSvDIxdHvcNnlBWYI0yRunWVC/1DAcV+G4uYTsSPPFawkJ56+
MNJCaywgCGPKoZ48K812NxMK5ryt0jsG+37KnLlx81MFyA9w4LV5mhQ9ggCwF0xi
2MBTraw4woe7gnz5Wwl1F/ILAJovWtPrvMdZ7R2KCi9G++zwNNVOy9971TAUN1NP
U0moFUdhsxKudDiOcss4EW3EAahiSa5WTq4DOqGYnhb1t3r+Xnd4QBLJRznXwI5A
zyO76a4O2HP6KTXrEEQaJFR3eBZJ75DV8t1P3kXbsdn/NIyrQu6PwqyAAPqMtvrH
HcNPBBZg21zAZhvGF7rsYaydmJaVzN4gkd579/F/KnfNVzogZ04SUg6V2MgAxUJT
mAI1L0bQiAHYPLmylnZFLbem+wc8RHcxfGQTow0wa68Cbr9SPyDtuzrPb+hw5dC/
r4tzuT6S6wNwfaBtBH/55lVm5x2pIIgOAZuW6Yiq8Xdrqq06g5WG/r2RlaUv00No
ONfQBQ0rfUh5D0L1C/mIfubgW2Qs+yGPf1mu5hpxf9IFoPHFeFd1xwPccT9SVHzz
qALxj81ndduFURRqoRocAQ2tj/VHvOdjI4Z+t4dva6+Sx/mxMVJolYNUoo+GM3ZB
1mJ06Fl5kyUOPnIt0zhpmjuHe3lSLJ43gDwEMnKdlPEiGiGXGH1h3Fhyg3YbV9JI
xKT0UJXkmPPbAXMimRik0xEXAJFRi0MGMPWwIYTyajseW0SoGuhfKl2x25QQ+iVX
WB5d/PiBCXLGEfOq0pGrJTboRFc1RsfPg357DANavmAc90DytR6L0Qg0jxQRbS+q
n97KUNFqEaMFZ5OE/3W7RdZFb/1hUXOpmCGRNdnpNpcXqzK1XBx3cpGdzxOp7R42
+tkK8kilfDruCjOoozCsOjrWK4G/OJG1I97zKC7ZB6lG6VtSvogJ6riGo+9z0hIc
ElsOH47BEy7S8LSDYrfXVPImx9U2hWV78sUcsVVa2c3iwneFE+xiUDposTH7qv3C
r5nukSh6BCkyqHn9X03g74D1sjuMHEC95i+4VpN4NaXS98EDD0HYgXig/aZyg9uT
B4a5Fz0bT3zAQzMeKUdCH1Y1YbSLqLMeyTD5UWQXa4HtY0iCNp6x3R9pg4FotcNX
kM64na/wBm3EU3+Wv1L0J/DxLmC+8uePrKTEVoLe2XF5iUqWvyegasg38DMSjMvB
0m9r6oHCbJL4fHZB/TW+wQmBgIpTbIbr7ucicTfen6MOY7C4rwzy+0iL3qE3O4OH
FamWya91tFzrLAMDvr62A49oSKwHpH7KXCm+q7hc/UMLnrCcWYSKOc2WCTM6KSid
d4fFoYmA2zVIFJX1iJ6Fy1lDu1lUAuSPGeke8VoLF8xtzmMB7sZBpm4XaqHhTIaa
MP1VujW08GuCd4hRDvjBijnoJjDHj+yuIFYzY0ppyYWAYE5xkZwGWqqRSg+MFYiA
tT7uHJuQWQ1/qsoG640sNlLAyKCwgr1Z4IrZLmI9BKxbCuOWOlGawmh5ZXk9KK/Z
tL75CR4cToQoijOWiYOmXGJMr7efgtxJL5hzVXiYOIlrgNqs4VkdmWqNJceqvV2s
SoWpVcKJjHaHc+mmhRO4iyIypANKq6S92NAaTUgOKE20rrWc+qNCBAhz65gyVoLy
zFIPOFwtDBsIUvT/2l5hMQizVt42dFDUtN4U1B3Z+TVwxZ1xq28xZhRzIFze+pP7
DC7SYbhfyOMfdCLcXn/vJ0wERd9oL+ixN0R2K37F9+jzNp4xJkCZzQINYmOtfRVK
yA1wkOJC6VaqMBZ4seT5i4Iw2mOddgFZ7k81Iam5RumDZ5ofvsCc2JcXf54c369R
uUv85+BTooNJ2vG9xOdez/JkhNvVcFk2hOVAylg8XD6426PdjvLGuoiwZezokzde
IJwVHe+Xlgu7XQisFG8asMvcipOSKVN+bzHZ0WU8HwUa1/OLK7obsdmtw4VwmOP+
kTv910XGJrgziQnCY5UwaOhQiEYBRkB5EUi//WI87w4ZDQDa4BTtKX3rMizaz+dj
SXDEWj7Xh2Df9NuKY07X97TLWLsWC7z5F7gR4OUlynrBNrL8y3YOj7nNyPl0aS56
1I6Vi2Ue596hmI48nvYNNU0heVyYUMAWeTz4rqAHFDccSvK1NXf2U18TkCTwfJoy
zHyvLiL4+pIXOK22mVWA0Q3xXXsGNRCsfnuHGKOzhUKC8AYeozl+Y42TsbS8PIrw
uqkm9dMSGjOayZ2tPZXW7NZUqDr7xhF72UAFWufgg92w5R0bUnsqLX25FVOg8mcd
QdMC2QscwmMRf7gObD+sfr1XzpEQUNV0fO5ws832LoIgwwurJifvpuK6tkLlgWWu
ucahbE0+XIXozm9m84eYS0AX2HWbyVwnde6QHQwoNFNF5qYJzG5hqgzLUxchDxpb
LcO4HvHrVRqvXgTCz0DKJyY8wyACDi2S8LBAItWvsd3LG1NSrf+BlehgxNyUDmyH
r9VCH4x0uNhcjeO+M1GBxkSiNAFkIyS9ozPu2/TA5z+xSU2zLfEeKKY/TT5cB0Ns
qLscZ/DpuYYXHIGFzXlVGfhImyzu4wfIrITV5D+qP2wvg6BEjYveH58SMRgMwaCx
vdbW6OmxoljHW37rUA4M4ow/NiHuLxGwi57YQhW9VoAvLp/0bQl7Gk67vX1+pI7X
mMP6oeyOD2PETA/8Jq2g5jmWkWzp+A5rfwTvBho+glHyaoY/ItP+SHYxJ3IW2u11
enesU/2Wje1XL1x9AIfCs8UgV1E4DKyLu8drquOX3U45zSTawX4zX9/dH1yT1nzI
b+m4bYQ3hHhfnjoOJ8s6Y6tL3BSzOXQRHmCx3Ftun57DTihNaKLUR56e6nVcfDip
Seklq5SP0oTjt5CscylvfRNKGIfxQ4WhB1Ex3r9ylNK8wCppnyoIsGIoHt6oviiu
I5tvSy5OF3ZNLrC6tWspJPsC1eD58NnxQlExMcVaOI3iCq1JKMhJ1tBmEwWKpqVL
ma6L9dcgkiNGZf9U1ajFtZTZQ4OJYfuhnvIT/gJUNDItSqi1K6TD/PBmbM55CmRa
3e2VvCw18TIdAHTn8y7pO3t/G+A9w3UTsJhnIVLuShzaEgZr7oOSgHXv8zZ5yaiN
am+hnfMqzUCzz98hsHjoDed0dnsS6kveQSmr4ID48vs0hTXvreuuZcINOoA1Mg0X
e7RbUt1QFsSnEwN4GDD/lXRK0Yeqx0iyKN5AQEh2pjeDpKKVx8XNIE6wkCk50wAg
pF6lbGjM6iz1uCb9gj7WdV+HhQiAS/VBLN+nQFptW0wgnGQk/7G4DZc9g6L6S/4C
bovpe59FrL9HFdLyvOWeC6YQmgEGyLfwjJq68oz8z1vyHCz5jEU9+qBG8hR4wea5
ecK06Um1Rq4ZxMIkdYOBzMFTMJQ0sUpZRUYr4AZPBQOEuz6EuFk5tctI5lzrcfzA
FNwvnZvF3j6lR4q6ysiH8uVIoYk11eKAxLFdkha20NEVSZeBDMz6RI3fO3fPApwc
SVir7KIf1UWH571Q9mug7RPG20rUXkXZ5vAkua5MjvyLgvjNm/baULky6W+mcNOk
IiFoifTYQGfBFuSOHM31rAId4A3G8BR6Hwt8O/hJ3+ozDcjxKbpnUiy3kG27eyik
F9Z+UCN6iAZXqZRJVqGdxKraC9mRpNny/q8BtfFGD6I4l3hYpHDBmOPd6whV0oYy
7DdJWq7NC24mhYaqA4LxV8rvC6tAfbBqXoEfLGxVwoa2bazTpzR0tOTqLa9LP208
z2IVbrJFaRHg81cGCtvpxUdaFvmkAv+myJ6buIzAllBZVxahGR76mdvVRN9LX4Fl
LR3yvaG3gAkvZ2/emJsA8H16XG990X7ZAwTnljRoAVx7vE8DldQt3zqhDpCuZxB2
pNHTK9gLv/pflmlLBW58JykCkXBzBxfJDPRTYt7XhenMWdTZ6LNWRSNZskTC6Wz2
I9co5NKbbh//5otZnfN30vprc/i/IWo+DypEf3RrOVdx+sqsvPXaegWshSpbVD8T
9YYzWdmT+VuT5wUtbM4yOrsULsyK5cXC0FmwJXs0NtSBYLrC3E64ug0OAouw47L/
uRV9+qRfk1rBDtukyr2aJK2S0jOudjw5KdhEtM8qtwqiNZm6nF8QErQRcqIFyYFq
u3yYDv8//mLHVGRtGNTGAqa2oWys38+/vyaDJBLjCGyEOmX/tomRg696s+34XOpa
1L9ZcMMFmAQSvG2HP+3QYs+pI+O4V98OUYlc6WeGCIM342sSbgqmfHc+BQ30S7Na
Wrgc3vG1+ZizdxjzPgpcxlJvQUVQbU7+Ou0xxqUClyQp/lyuJQK8/uToq8GoZ6AI
AGhRd4rz6toUwF+cbJ+gcgez4+v24YDkS7QErBTzA39rT3p+f42hTvCNmJ91qC7E
QZdquz0DmIKclfBv5zZGYXzuvWWx/MLUSnEceLBRjF9H4KowA5Ete5WVDezQbs0o
Tg149D3zJhihvVvRSL/hu/ODlsgI87GqJXxvn1o9CttSwJwPywZf1wmQ1F4IMmge
dPhos6umcyhF7cyVAVX1uElIA+OWFCTZV5ssQMLWNqicG8+7Jcrvseoa/OhusKCQ
c7cRsZKbvajyHrJ50qrg7jdVOYh7Fi1nFC+9KjAExEXZ4bnDra7CfJGs1mTgFElu
gZCYTux3fk/4YLoa3Df7V0eEtHREZ+J7zg82inCbBhl/ZKecMHFu9YAZTYKk5myW
TrGV7gw5FIlQF+CmwWmjpSetEOVDH2uqiZmFO5C492FKqgJF6+BBsDo/glZpFcXv
wmvmBgTu14h3djzQNjCdBO0ewEj4f7ktT1H/NXneWXIlLxixH/575um4uJMDX3mV
ncwWxPu6U6mvNIY/NQtJlo00VpFTiwL0qH/xWfLey4obNac19KQX3oTt0eHnINog
bzI939Dxdtwdj9AvJzKkqp7a7zK/eZGf7YWgMeP3QrPg+Z08ENl+rpOeCmx7cKyI
CYQGnTVDxV2Pu+mR/KigHL/HAtx2HnZIA5Hc+GjpJnD2uBJdCzD7N7ARXE4Uc0Kv
I1PppQvygAq9n+wZpfkLxbrzwsDjQiwiV7sPhIxu7FySWu27KyMSDTq93IHyRbeU
+Bm+OXH2Ze7Pv7qp829H4L04YqBPsNvvvB66SWE5KeNsjOuVJeCJ3T3bTtDF29vB
alQAu6Vauczild9HamVU4d2HGllWd0rUuurjNqtpshrvs0UnrlG3tIHWstUD93h3
E4x4VsXwiIAZot+in9tByXbjN1VG4FYDY/Bym9C0QdKTaYmomxNscaqeF1A41/v+
c4ZRZyY95AJst0W0F8nxQZ+uf1uuLcen1FkYR3NGuZXEQKFndsNOXcU2bHPI1UyZ
1UhsyUxdiKSuAfCO0HDV2eM2cjOEBwc7ZHqYkdPg7B3kM4D3jdW0NZiS5pec2ihf
1F4g9/vTs/zf93mWeFClaQ7P0HssjTusi0MJ8OtGbTd20ZYUMdHMJEViJwmTnAfl
ukfhpYUdnEtBOHvdeCWIyzNtNbnN2AgaR/qlwE50zHpvoDiGR1qCHkQULHzEjSwV
PqwIB1UGomr6C1nQH5kpCTx4lBBMr9FUrKMOOJ0PZef9Iaq0OiJdE4DAIg9vcos+
DxUM1RjHZlSgUTO+rgFOACwfNW/2KP2AHXPtHpvHHRvX6xXudShRJ6cPDrGiJlY/
IjUh/w9ANNH9mXGF3Isnqb4Zo1iQPdivOUZIkoE5PvzNmYq3VUr2P9+duK34bOAV
GGmmumfvb828KZZaMdAHYteP5cowUlw8/IG2mHLhZHZASVKMtDehSVsdaieitzDS
TiTA47Ca40gwUn00XC6//gGnL7qy2rXOYtNomOwoaet01E0ju1gJRinDYSaRvVbO
N46q/FwQ8JOvZxsSzoBhlf5HM1jZMf/Mpplm9WCnW0ZhmwsWPWOlBLJwOddiS5gP
f7V/dd14P3x/KVSF+RF9zNwGGrvzZcoENB2Fs2Vv6cSnV0bQx9QRkVbJMebM5Opr
ra64CmDOuYK8FjegeYp62ABZiFku7G+ubfBfSn6THjm0Ieg5YwD4Ag46QbtQJe1B
PmzzQ8iRopp6yyI/Qr0oC0n54p/tPqKcnXthmP8FZnwbA1+40lJMWS/5QKDerly3
B3HesTGWcMWw9zVBNHJHmwyObN/vQK4/4NoztM8v2I/7YEcT23FrUNbPVxuo98DL
oWhJZ3ebO+V6LHJTSiaV6i2Sj7/wbynmpqBrvvb7o2PBeIGAy4Gq3qsH83IfEY3S
J55cdxOeWQBRHuGxSyY2fXmn2urgGza6gqvqkOcpNurCPh0dH/9RKiP5VnoDn6D3
xYIbdupsm9+ZUlyRkVh8EPeBq18RBgMxf7LmPNQkz6K5ThAZCrGFaBXNZFhwyhX7
5h83IAMtf13plnPDdWWKWyR64vugvbdhmE/SPdL/Q/p5j+ejXrbgiHAL8RmQkib2
MWnNioRynp5XLHuSWQOqOuOZyZ0W7CE+/V+PaNaz8vscsoi/EyJHvOJfDP816LC8
JxOBmp/UK7zUsDVilQOtmydAqR5wVZu7snShGI4QfFyz+S6Amjl+EUWZtkSraUur
lPUSlcvkZIgu0T+rKtqhCCx2TFBwDz1vvLAf8qcAbZrmDblQeifAaC8E8Xn8SODH
zv2zNpb26R+S68kxPQ6CT1B3q2elL3dZubXtrjJUfiKHENubzi3TzFrhVaM2UwYg
uA0OqnxZHPMiVdsrVT5h2/uxvGVoWXw0Z5ocIKzT1j0qk9Zb9CIW/tiInXENevHY
uiYoGI6+60nq0jGmKdMCZPc61vQDl+GUUEtN3rfvayvSSelCOk2jw/EVNnsD88uD
Y5eKCNIWfbpS7CsY2PalwVMD2upVdFC2DAbf+bT379wBVfCFzK4oLAwye6oYv0aT
mtV6JnMplkzMo5sAfL9Ui5qb8ENGAoGNtxhvl9uD2dqHnIdPiQblp1Ddbxh87Wto
Ihsxn8dxh0pRXrA/lJBPHKbT0HERXyVxMbh1sS79pMihWdG3NiyKrK/+bnaLixNs
fTbR9sxXQ102dTe7J0hGvRkW/rREt32pPPtpCGo8nXBs6MqBmUdCYChGXxtdA6HF
XsyimML5qbe/2EBGdp++jTNe0eVjs1iRhqbV8qtd0SPnDX7HcPc04fk+VwFPQSXv
/OhTbynD0eg2KO+JxanThtZMq8xGT3hY5Kf7hWcj7HQXZvTAKwyrOgdaFzuogU2Y
s/95kg64WUlsjSknJp93SzHLEueJf7mqPJnjK721dTxFhECUmwn7OpgUckUMqgHg
Hb9VvC7+4pbJ6sTooIsbE7KKV4vBRv7V8sFJFBWh67uBj5ao3i6vZgcFNkOsSgp/
9WbNs3ttVDH4OwWylRbqDwbAxKmmIkcPlq5oBVQBkJBmZJs13XVaaGKVfaLaWLlL
dUdEe1uRqtJ13yrY6GqyRt7CPzNde/UWlBV0V7/poI0HrN5TyQkmjK+KX5Ez4eBd
m5jHASsHGYOhfdrVHfTZN4xwoBlhmwKeNkR5bO5Q+7UICQRH53bRuixUI6VH8zxc
0ys1puk/kw/AeJjPBXSi4zkVtJ38PbCiflHi+Q5D7lvr8LfheS2/95ms1JtEAd87
2PxITro5v1jSZfqQCiXasYLMhPwaHtVAiyZnM6oRbTTdwbi7HOedQd1G3gOYfzIs
CMorkMCjx+/kWHn6kkGFv2LN2gVGC7KUcj8Y4CVZ+T6LyRU/y3imSo2cpI8HK6b5
GWGcEDEML4SCH/x2PgSJnlP7phl75jRQqNMOpN0ZTf9Sd4CDT8q/8pW/B35BWm5E
RUV/qrsAg9DY5uve5VW/m+D1/EVorTrJDLsYJjcAwWjigX94X2aex8J1mJmfPbNn
MkImph3n6H/btrEMtAVDm3ZjLai/c+NdycXzGrky69ysWptocgPdD4xQV8f/Tmfe
3IRRwfkMkuFFh99Z9EhBsoS3RUjK/4jdek0v9Hs8EdnkoL7IbsHXPdqp1jgKovbu
w9IcG5nJZJ/ppYGRhTh3Z9myQ4M/vgb+YiHQ+Y/QebIp4paZjkKvUU08E1KycCMI
nzpX09AnLKJiEWC2blhEOyTwE7LeHFSw1RusxVwfTO6/OaWBxcKENLiHUu0ctd6k
PYbADpYVbF4Xjek6sPV/jvNpaFh1TgIp18r33m2uqeeKV3bUpoREcVzUP8HU/56o
VzQ/9YOTca5VkhB4JHm41AAUjvAAZZV/SSdypYyb08Ma76f1qw/fcGOvMYLdysaI
xTuimaCWJRLJ07lCD6+V/UdqKhKgu+Vh0wZQGhiyfUZMtqdm+D7eUtCJah7xCZMO
alekY0wnzFhrxHyW/BfFJwxwElV+Xfe7AHBdYuVRCxBPxQF0CpXMDMYjVesKbH99
PPDqvjy6ctR8Ws/WrsZ317zUcitBXMhz+yo7BHVyrSLwOKWCxe1GaDmZtg9cl3kl
0meJoCglXf6XYf+pzLwWf+MaKj06Jd8adtInwN0LF2zoflC/1j7YeM5wcaEpriF4
FLevJA4pKdkDJe/4plzjoc8XdGCO9praHTLeNx5wYHwqFLprRguePOyOpnoBOUP6
ZQxNjg4sA32SGmsqTF9dIkm0GZAjcq4izRpA9B0cStv+J4ae820sUuK2R4Oj0hQt
0+Kt4Ez8jqVKrtlYFNccAG19A48eOo8RyQp+bk/lKZ9hzGNqCwe/FdAULC1OymR7
ZBSb37FvpYlyL/BnQd1lNL8AX+s7Hb7xluFvnuBWUdCE+J6nKbVHO4Fbdu89FmE2
D5wkwcYP2a5SR6rnLng62+UiZLPoFpjxa97XW6nPaV2uQ4yLKsTJDnpnNpSt1SA+
FXoDRtaONLpBdo32ESYaAZUI7c1LpTNkHw/XjUwOppPp2Dk96TVNTsN4B4euJS0r
GHPy8S8kZC8QEU6qb/GpYSIhR2wN9/AFcGLBP3N1HHawJaFeXm6JWips+3VYasJy
f1ZoaSWR0wogkg8mG+RpBHf+Otf357jwJm3Siy/zPVGcvdcEfRYAzhzZDFuEyjxy
fAOnD8ToLDwWUQxR43LM1P4lGKmBm/xiNJ9yEJYlbmpeq5WojD3f+RGd6AI36EeY
SQCG9QPFIYFwtg8b8mQ8LfniltLSncuNn6VclMA2hL57yZDgg8wrW25tZBZxw1/S
X3D8+gTTDGsZDQiRLo/xx79DG0ilwVUSjU3ulXqh37Di6WINZ/EsCmNC2Xlc9693
L7TGcbAPiMVbSapQ/8fm5hOHg35nCYle+4NE8MSAPGFdGM/LoKbzThmlN+d163Cy
lCzSCEd0AJPgobVbuQbEfeB0pyohQLXbyg4RGO53HiU5DCijJQT5Xgp6NU72o/Tt
dvy75xGSmiWAAJLFazqQMhG8/tv0Vpi2PcRvsXsQE5bqMqK0iPw3+BwfPweK438L
ZYZ36kc474XuvrVJBOXLtG0R7Cd8fX9p5AXjcJv/Ft/CkVNgcOrqxqOTatf7W75p
Q81IT5BMiAenrI8lrKIvhaWstlvFrgbWqxxjVJvHiO/EZzD/VCeGsH+A8hDITXwj
ccNAPt4yn1SjXW/WBZN4xaYOA7t8SL/dFIVGC8EtoRVNPWRpCU8foaRbnqFhPAhj
zKGgb240/B7C47g3KMQiU198GqQluLX9DjCCTkpIq1WP21VPa2cs5DmZj4K8aJ9Q
qlGdf+YCYGAMeC0UTQzOysL9NPm9wLlEsLY+jYwFpwP9wq1ufbUWFzCAZX6U0/uv
nDklPpHPQSKoGPq+nh8RnoyO9p16dEqJBd2mi1oITbvGPTOEyQ0SDMaTJ0JLDSAc
T7xYgtfP4XfB13W5JYMvrHO/7i+STwoa3L3XWggWtEK4Qt10hac3XcjeI0Ss9Gj8
H4BipgKvq8soYWwT9ge7pNWZskIs97utfJfmeOOZK40YeOv54lz5RvO/eMf9eb9+
NuKdh1b7PQs2c5Pu+xHYm3AseRzUuuxNPySBBIa0ilS35qVZi1HHGaO7VNAGo1nG
lGnIHbpHphzmDgm5gwV0G8UqJdFj8mLTaq1zTG45UiMGj9JgvbJmnbznjgeEKs3r
3FA2lzMQsR+KRPeCQdFFQo1IYxtajv0XNmWRcJcIGe9zY0WvFx357+Lps3cgwTdc
sc42Jfat2yL5dlQBzYHs0Bef3vdLGeBUqFyPErTIrUWQSkS2UPfwCTh9gOTqu+f1
DrqqMqg3clBZyKe8EH4dSg9Fq2ZGXqElsW6Si5Egf+JO6M2YjAE+Dh4nlrxaZqha
SH0S10VVMs2mpHM8zl3EcQL3rgOMcAQUXmzKFCv7snHhUefhc9lf5OJscd0VVY/l
ctwTtYB11TaKyrhxMuJtrNLoNq9slMRu9YZgMXfapiZO1Ozw+O5TA7OmYlQcvKxQ
jjgPRBfghNqFaH/wZ7ULgmDmZBHC7oW2HSYwoJpNHMAzwflGOKD/efiGm7+QTWyL
PYUfm842k3i4CzLBRgoT8TMzjxS+wYnyWRCl8jeLq5QDsBSQ+v8hNIbqT8VJH7Ak
Zn0tRKkJIv33KCeY5vHiX8Nz2jwqoCiBmDE5p99SOS2CcbTW9z14lKBS3iyQ78OI
Njg7M2p+xxiBv5tHXpJFK91vtosi7Q/eK0OEVe2fDdWnLlYc7JmqZ3x3hxH55YlA
Pmhq9Yi2AMDP/ZMhcTMXFjoo1WTUJtF0oj16MSVQ7c/GAuApBgZ/XsIcCLs9IcKU
2pETqwC08+Zq2Jil4dyoNBOtfkJcf7Vlmcs55ALKPunr5EMlLawR6RXFftDfdVMG
u5OfbqpHDn2QgncbmpiQmszoGQXKZDjl5+ZnIbPwfsL4W6sEbwR15j19BqTq7jdr
LEQ5HZ+QPexdMuPm61RUElpdyv7xWozXYl4fN96IcOkV2PLvBVqLZMSMCMY5h4B6
Bj7JaiMwj/RmQvrNygysbJjEWK6qrkKkLy5r4Liy1RwSdSrwAzOimblYfsWjEy+f
MAI6nnSk/Knj/pApf43//x1voj7hRFTvXvOAYA6jE1dVpS9f0Bjx2grSc6wZwd80
u4GTfgk62B/g1RpXkcMeFehDBQMH91UnqrZNXnM21WSucirRaqLWEamN8SUlLytx
bH/zoCpWJqpb/KdzcEBSOIco3BkIOo0IV/Ph6VwOc2UI//QKsTcIgkOndRexi0e/
PayCfm8ZC08AEvgljI9VG7HotxEL11Yk5FeI0FIf5kE9h3elQ0zZe8czVr8A7cuL
LtZeIGP3hDGpFqzQYPgBIiVvCwwr+z5OIPrmDT0y5zs2qzjOQ5LXagVIRJ3VMi0R
qdntD9bBij4OAm8kc49uc7IfGWs88VnuoDw0fDBjCNnDWuTnu/wNltpQGMRDqWdR
ZFdLiWN9FFLRkH6ybq96tJO8jy63QibuUYxQz08tggCMwNyF/bKKkiccAiC/z3Cb
TIDS7WaLzk3cKdCodza5WzxR4aO3kcVRpjQ6fQhNv129ng/mKf9Gq1mfWeXZbsVc
2tjJPyT9UUbIAleIsD3+sW+15Pkywoe6Ysv9m3uvthx++6OqFYGgZnWINOder7F3
DzvDjNKMsmcrE4rZGTUATC9Y3lUO2HakgnNZzL8d/kkR+jk1/zjl0TQsMEmdEN7l
gWb/W7zIT4464gx/CvT0duAv1SMK0FOajRlqeYB4qI1r7Qk0/c5JsvB5+CdWOzyl
4ZtL0+dJIz0Q2E9kHg48pbQH1c/PuPrUhDPQoKFJhLSuCg9fh3TNOsqTUtbvoXbn
V7TpsrEGzU+50YFRRWHHlnleQ1m+VS04GVE5B+SppGLZYK/ICeW5B0fNRSU+ROvW
UzAOWl91ucGjGEAnEnGKdDfMyDuaF5O9ZQfTEGDO8zPQhsPsHp2Hm+nPYVkvrrOb
x7uOopP+Iykavt5j0/L63F8Ak/fGmMdKq348WdUgQ3N3BR2rnA49elIBJgzafnsu
Suzs9Wx2dFlr2jkv9C+ePsgflQ0ZEvc1SEVjyHZxIYqugs6csu5tZMSf98DVB/Fm
ckVk9VbEK/w2MvhGnIRl4+t6Lql7rTXaYqmh/TvhfcqA0ZvjJFOgEIZ6YgS/gTQP
1V2raRXl5jDrYC1ouTr/g4hNGTixvFJDFx4y8dAOUGRrGenTDePQXfwoPpRuiZKs
TYOPneMzhOWd/8SOUwdmfQHT3EULE2DM/2hxhBQS2oRTkMfLrKJVvEfA2NH6zf9v
9G89k+KXmCBn9Qus8gHC2IJa4ML3PH4sX5F22gDDzmonoip7gjknjTIJ0ZKj6TIK
k6SaXT9GFATdCUk5BaOXBhONnU0xOiqhpYMsHgoB0JD4+yghqlrxCw4kmoeFoykM
EPQZyOfG1yCgysmaVZ1J0q98KowuepNLUA/K+5Xz7KEu7gx+tupvWnCiteFr0ggE
/FgvdtHyLv51xXI0brX+BuWGQ1/tFaDLEoJteBQsa3JYPGT/FKJXTBvyXlGbQ1AP
E8OFGy7kRLVZYvBOa9t66LXP7XlD+yw8v/2weSfvjjTMHUoRhGyCal3AMde8h4LD
U/yFATDrZ7gtWvE4iOPmMvybCpunnsw7rc85QzPXM/LpMm5jliZLsbCajaGjx3Xc
ViTcFjgUP3ukt7eJtBXcgWj9a7MyONUdkmgLscnHt4eysNnAP1JaNqrKU17VJjAP
zyikQHzpY873LOJlVlu7kDiAdmWQUXprNCcowoGYc5YBP5+5RPrlPnJO1sPK/NQ5
HRDGNu3C7Xy6Ucq5JKmArDowO9ZTu5RAWkt74O3/PlirWy474rxoIaQivg8EkZsU
XIaWby55FbUnnVi+EZPJb66NI636swlqfQL6PpS5Jc4UUWqHBRXcFjBAtfhKFSga
jmxbPhnZuJ2ZYfq+hZAJMCqTJvbbdgjCG2EcFVgBPv9kORF4MAKL6FiUOhXf/F+4
cfO3ZgaJzvRpJkODUwjqtQ76PdjssiBgkswDdo1lrKSqwLv2YLU299E1iGyYkmS8
6FlBYwZzAyshq7pEMMbDbLN+aDYZDp75iCM4akO3n2hwMYQtCik0/hXpxCXVYVDh
zXTKNHNsluXeRawqIWyfV1nW75L4QAOnhir86vT08sijmCZw0f7GQc66cS+/w32c
MoT6/l/q2aWUTmxMd18hJrObwsMsg9VgUPMBHemyBi1qNoHpqlHSkB1ZoHa5YOVn
6j78XDRB/uCkfDlvXzja+m/TG719+/Xgk8c/R9D6MFrcCHhsMi64/uQNIjcjNKph
20bkjAkPKw8pZ1C9BzvGdqqOdH00BEvHwczwAdFO6FLrZA/hPt1MsJtt+1Q5RwDu
doOgmcmL3jHscUmb3XQvji+2RSuCpv+gnnUKJgyuNh09enVzshBY3A/cqWw9S5hI
xu5oGFAigIK33DY+CBa08eU2dfmt6LzrmlDda55Ku+zOmhieI3TRcbqukXMxvC+P
k4/YEvZHRk0/mY5r/LsBOEZk1vkSpicxr/2CAZ/ArIm69MjZXnih+Nn564kU8+d3
8qgrQUlsIhg3hP9G0KXjqSKxhMMETEjc8h+b+QGMTXdBscneTsVCpeEVcQXA6H2r
kcg6ALm4wn/hm0WXsKAmgZTXzhPVNyEmM1OS4UFEFFPZtSWTTmDr7/CDdErxFAcX
Lo2quPo+Vg/k92SvJSZQOqaJIvJ30jDWSYZf6NYMYV+PIaln0DZqm8cOa7ViSLYJ
kPdQbKF+AUI539aolE09L7HhI1PXrjidyks4CXN09uBQBGHeNPyqxmj7ROldSmfQ
wfp9CtZ/kTi232SBjda2uQdK0/rVvQpKGSM8jgbNMfO2u/n7i/x79BrgyHjGNY+T
VpCVKxFTo/bk929ZYMxpikNCq8nafJwKfZgJikYxTQtQ8ucr0vGLG7AqaB6bZdsh
DxZs4rhXgGJx3dMg0UqepeWbzwbWAB73zYZibB+b/IsA5rHZMc/N0GllXc0xPsMA
hh1SKa4nYXjYutXWh1CY7DT+yZruQl4F552emeRDst0wOtSmrCZhu2YS4wy2XfG9
qWRKACJHOM4fFLsHnxA1xmdXUmZVC1xH9TZ6CAZvNHFrQnzlpb0HlSugpz8WTIxR
kRoCSeI76VnEuN74UHjCxddF+TTbXeFdZWQ4IlXm1AyR1P8T2/LBk76AVlNIP3Et
JkS2MtUoDsh7Ojtytisdb67XCEoB96KSAQSx+Hmq7QuduivM4c1nr7Kj4u73396i
wSTo19xMy6IBVWaVwgbaQI3qcxYLU0slV9JMFA2nJ1bQlnplsLkWArKXZdF8lQhg
KK9roqNVQuMtuhkut3uEtt+2HzeuRmv4uTZlzjx9jLDt7XSpQHcpYGbnOYxeGsbc
ZVCloGEf1FWTgfptFu9eaLZmT2Trj160U/+Cr9OyWks9vbJjO6BylZaPZp23SBMO
Yk7P2nKhE9Uf930P4DuH5u7eSvU3gFoUlweonCGsoRj8EzlfcglA5HM81bP3Xl+Z
NKEzaMBBr7McOzsugyFoa8CW3U9CP5m5dv0Dk7zrJcgjQh5y9BGeoE249VrWZP1k
Ft4b7bIrxUoLpC2/IsVDe/FZbWKNAgPkVRfmFtQHmhz/f/1bd2kaKvdLqDZf68RU
Mg9rnuqsOPZGJm7KQkRb+Ee0GtUdOSkTmCfy1NZMRu8i+UxpGWxLQ3vk+gOi0qMz
PgcUrY41OUHdd8yMnkfc8o0hPTm/M6CmRyY/YvJhiB2bUgkXh6PMpTyX5qFkEjij
bDRnTrX9CRYB1MrclADFgoE4JH4Myugm6gp6Ip/BKPZuvAdOlUuSCPySVtNcTlL3
pSaumUWEnADw4jcXWavUgzGxdp5NDPHosmunIjlK/D0ucVcfJerU3IqM3bZdBiEW
iG+VMulLdtQ9WlT7FIZdCw7615dP0nQgR61UJTsSpi4MsaUkIOqAI7+ALiPk4Ijx
wfNOs2eCsmcmCE1SLWWKpPFBIw19PPq9AeZZp3eOd5FPAQAqWhVrwYROFjd/4YHD
3Gvtdi0o6qyD4jMDuUyidFHlbh5+9DdvrT7sXdg0wtz26PVGs3Kb8VQToG8hCC+h
FqG6l+MfH4XBS4CkHvQVH5uS4Fvsshsa+y3D4gSAZ00KnaoWM3wco76VlFMDf5gt
ZmkqXjgPIRrzloO3C/3vyzv50d9jTg3EX+seWdrFwzAXCE+0RcJkhFdwqMTZfC/m
g7toKS+j8/vjoQjuA8NsvEEeGm6eJPVm1dEPgZ5+i7iJXtpz2VGu5Ag8dhdEvEdg
H1aia2DFGPcw0T+wr/cw5Ehv65jJ8ELI+vvP9Jcp02z/FavakG/xE0u8zMm3vKrf
mten5FNXU2617jUjcUK8Ua9/YY0DFw8b+JqpHOrnJKRDwPmhYXjR67R7Ux0MBGQl
kk+PT1zBRn1d/Ccv9yYU6Mgn+mc9UXjRTKBAR/ssIsEntn2CzDY55hnu5Her+1E0
45sAVOhgnw2kiqsdaYrbNrsWh2Ee1Qs1JlQGiOaKh3C3vdbqxWWcXgjkClbNfImp
JIU7vFxi3fwERidWXpR1CnYPZmYAFdq45j+rJnt2YPMGG/JdGrjd9Ax6F3enhD9+
MXmYG6Lm9LlGYTsMD6ebBJuVasTbbBaj2Irfq57IBqIElia+EyXiYyjRynvn6tNg
iHGImaMT3JJJF0YB63pCAaOl/qsZ40wlXwID35UdUmzfzSYL8iZ8/0Zl+2s5TDZc
2GA0CJsQ6RU+BRNlbu2ECOBzrGA+YVRBR0Ri/d0YsUmZFn6ugVY8F2g2EN1qpkVe
eakYWHA038MGe/m+IWwGKCblFDlnjScKxA9DjWonErEEWmBi+zWkBpO1Q96EdTSG
+y6SpNfP+qQseprrEgmZV0RCg/VGZcTPyqifkswzZG/fEGjyhWp8YAocr/dmoFEJ
1J0c/yYvokwGpoibLyzcr25B5orZ2V3hy+bNvhC8C4r/olWn+WbJP1TWioDjUypO
eI2KaRpwhNrEREvrk0Te3pIbUwOopWL0Iet6k4NRTULgKezAH69JKpiWdbvSb94t
G5hyo0Mc1ZEdkKDtraFeV/zsHOX/hU+Arf30MFa3ZJLL/ieku0As0cvKLJb+C1T4
8vVmHklWj1s8+MLxiy5nNEyA+xt7C/Ds3n4ZhcAm5YrWU17/hu5yb06sIzf+xNe8
KcMB633veFNcHC8ZnJaki+W09BZP0aXyukkW3xRenxAxo+b5FRiHpwa9fVi5SGzC
AHt0pooqiB58fHIrK9PPW5iCiYEc2JQyKcAGWlyrozfpTwGL0xcft8Yfu2hNvp7U
41D+xFvctYuN6ZYdBLf7xqYUAHvCWVYLbV2MC1oScdU/4+z634QnjjOwasK0gHAr
3pPLGoCNgT46WGWcKSO9iK/Iv4ppqGd1YPUW9cUPi5oeLLzFT2GtgLd842jbeeGM
PgLRr9D5iXE2V2oefV7JpU0PRDyA3TMP6gc8xB5O5KkK8psneDlHuJsnBQhXntip
EVPa9Xw7lVPLH3LUSrJ8zoarv9i4XCcnIu6p5nTKtVVpSJStI2l52gxsqCqVdLjs
wjWLr4p5pLDyroQz+tSokvqU5yrCMgCv6yyCXeEl02zsiE1G8Q+Uk3Gm5lbZwrLU
H3LIdOn8lnY5WTEZCdfKi5c3rzq/9qFbYzGp7f91bIoGjN0k4jDyo3DfC07CSz6k
Rktil3dKBSoJVUPXppt58wuJGhOrZ7M/mPD3Aut03Il/Lf3jcZNu9qIwoRcXWWN+
K049q3eou1SLPhe0pbwkALxfaoTz+GOhSnLfkCoBmpLD6PDaJh7di7GDaZtVdwdN
22spI6Fhei86Pcr7x190T6e+MLccdf6zUAH2pDqSyd9HCwNxORMYmhL/Brqo9i9P
YoP09jua58ZD6Lsb/QRX77236LzU7aCKLFFwk8+M/22R/awFp8LrZnv2TSWrO8YB
h+Qqe8+yM5aqO7YYiRZRdExNQv4oxNaLupgDT6S2S4RulpCMYpPFNwC84IgPROny
05C/5URKGbBdrwJLldaw+35lJ6peX06kCL3JTGbn4cPcZh3AYcaBoyFyD4jMoAzf
Oz5PVltLvbBheiK92L7HBplZecRcHxZz7eJShjqpbxNa2h78K7Zz5vCloFuqMgK2
5/CHIcPTwgNtnGtej0E/LeNVale62u+Sxfw7EvgaIQOxkDQ1bVVhZ9vTkCdeTDtm
EQ68plsazyglj3r4fFEdmEI/iY2n6yADygl9/eVwn0rlfM1G5ZKDCpRkEkCCJpAe
34r/OcgvNsDFVbdi8wESXNCek5a9j8cGTmx+ig3NFP6sZvAx0LtFx3rqkd49lg9W
meCgLsQilIGHdy7s9UcGpuYx9fqW7jYE5+41VXAgZTE6VS1PK7jeQVly6ufHW1c0
GV4W7/y9kJ1siSHTh1l8LVNxnw6STxhviCfT3NtJdwx5IBDHOPBsMefQ4p8GvwrJ
QHhFcPhBMrcu95wPX9I641TCtSeZvRLoLlTl7L/AGnmvCh9qY78Dt5cFQmGvbwn3
6Ka3/eV28ffJKjawJ4JQNhI0K5Y6qpUhMA9vhDOWLRsVSZLwOqmSRbeetKB8mLGV
+qfmzsLtZnWsAtn9UPl6H+RE2G4ZMl4aYkVkQtEenCGEiHTnIKm94PTObrr3mbDf
IrR0ENuB4KBHCq0fGGjz0myCufx1weNUrVujt4OJXemaCqMT2aROsY0IFVtyhWYQ
a3XgOltc/5JdjAoIiwDxRbigUKmQCKXz8gxQbuFPYy5NC8RzdGGj+Id2SHxBvSRw
xuA8ExLoguDzl7KWsgAYj8DbvjgMS+J1A3Jf8vVY/AJ8KRRg9V+wYe5nYUkwWfCk
mMiNiJdRF40bZC1f4jCrUTqSPdCG8dekLayl9kg2C3h1RgXF7RpkPkGV7J106grt
OTHAyonshgZmSJ5619vez2xwfEcMjuo+EAMhhRw4h0xP+B7ZF8P/LyVZ2PycWJ0M
6zbdGdCSQ8XjJ390jNAXotdkmDbZrw7DCI5y84nYWLK7MxutMWq+7ZvpT6Poc2jP
GdKepy/gqV6QdM4RifAW2wbOsSoDy+aUCRlukTi+5RXavHMnMEACEgtLTmSm6Gwp
BANaUDE5C/C+0N3jubUOTCBa/FnkLsHi8YxFhPcbncWVFUNq8TtiOLkbmKW0cOP2
a4Q6K95poZNobLXfbkHIe4TRREyATzriXqPmwyvBaW/weG5lmTV9NsYvGKfgzT9E
o1RUsndv0UNmcOk6oH0NfVYdetkRiUwBQxUlLpcIxi+cwH9tvYG6HvtP23I5uKxo
rlAZbLMHpmZdPoJ2GZFAi/H8rzoysWznfz8jIVB+5rNM+LHvKYTdEtqo5FHzZunK
evGBqhJvKMiYO7lRSF54tO3EtHpDHZIYseK7B03bCeWgt5pnkXUB1Mq5efGTrMJh
NYp81NpvfkmhJmXgNeAgi2uN9RDMB0OkDB7lS5OgCURfYBYcjvBt5qZL1p6VbCRh
njZFTzG7429T+Pe4C1lLbwdbw44xNuG5dr20dGMmkHBUZ73SNgUJgYMHwZ9b9X7x
hhvykHu98IsA+1lsa0dAnJ/esjtI/kUtecNoUa54cAC7BixEb74Xf0W1idub4oFn
38Sumz5vbYPNLqSUiL1BIdIHNUis4q9hzvJFmtNu3jtsF9phuanEAGOsnsU9wRGL
RuN9eoTrl+f0+aAqYi0JNt7aOjYl1v/EwER9igjbPjHR2ohrpAqDK6GktoY8Eku7
qre1BfHjUiZ9TUgTJXj/cjCb9T0zWvAdsnaRp8nybTifoLEy2OItrjwDZRMQguqC
mFppoZeUv2yFcDQWMKjJvNPcIEJfdIGFjsr9uKJbKkK1Ig6/W6Pf2qovW5nzCOBb
Lpua0P34wxnzMe3QXkNaXBvk2odeV1qOSkKSkuDEYf3h4LeGLKgPDG/Pf85Ec9o9
CcIG8R8ar95Q9TzJD9+TTqmLn7/2OrnRtq77F34WqmpwkqbXBHHOrgqIg54PVKfp
hDGW7fpfXIiAhgSP+8wkaoMOLR7Xf6P3imbeZqpTvy8+k0ZGbKYtpqEkbkVbyn/F
jDPRLVBzgpcjHsUOR5BN3Q0tutRqreZ+tc0tAiBUCp591ZSXta41lXqmeoIyEN41
IpuJ/w8fSAsFnxAvDkL9hfifW7UAxL1KQjuASGMy08hfECbqb+/d8Cl+w+6WzU5n
unos7ixtAd058HS7IBOIPjIpOgQQj3HnWH6wSZEZGSYiapFfgBmSumrie+Yz2Ii3
yluB0hcZ0oH/tFh8wHVRhDH2uuCMvX3wcHacBMPOHFqFChCvJGXx/7QJz79jgxBh
Gr9Oqq8fakJkjefff4s2Oh1g8itvhhzGG9etju6qeSMBuSj6zKyZ2OtfwH9TLjSL
76gHX4pJ6jZBqZOWaO03TcxEu5az5OUjUxxIs7A4IHsLMxioWq6QzmaQHqsMrtFk
KD7hxgCBPt19R/KbvZK/ergwgiIQiQySgZ3278gP9merwBQC5yeHpINrfO8BenoN
wg9OEQHS9RyQzl7xFaB1YkYBMq0PI5LAu2QYpLsnhDnILBjce2x/uOqR4cfduRCj
a6sw4mnhFFPEU5YYF20fGFzZOA2zoZQxN6jaUtw/48uCb1LQaNp9gSjoDG0oeivz
0uMRWTA5ntkgthXy38sZ0vaZ9dS3JShuX3ynMZ+R0qhu/zV8fySD2BJKbGy3veFN
vNjANbfjz9NlmYkz29TqpbyJgDJVtEoreKDyd5qcOCaJI1AbK6vzpNc+rAEWSr69
zjrskRezLIpoCuQKHNpVbL+qhH0xEDsGUTfab84JQgRBbzIxBn5nqt8ZuMZbu81K
NIQDFC3dsSVfKZeaZ5NzHosnSLuQKoMWqMdWBmVk9dazK3aPhCeaZy487+zJOTHw
Z3ZmSEf3nhvfR3Lk2GBoaiuhshr//VOPTRx1Uc8a8Ld1K0Z6eFy85eey3U+EUZsp
YUhzsiTXBL/SCtml2sLdip0wL+A3wlmHfSITmBsQcQz9FcvlujPtTVjJyvPApN2Q
uW2JfMAxpdZ2pXA9UjRk9Qf8tuWJuKoILlE66B8G1/8FinV5moll+okVpSfkjTw/
gmLEwJY8OTUnNc9Av6aZjzoZl06dFyvzrjMeCOONCOcbwzw+zeJe5w0niVdEn0H/
9ZMs2k5IlTXnSbJdUcrZ9zM4x8JG34hOk2VdEwsy2+Hs2cjHvnK7+qh3XUtVSV00
gVyK1dz4+EZeIIhkShvZYYueDYY5Dob5Qyh0OTOv+Mw8iZAfz3SpGvFoqIGKuCoe
MVuNOku5JRpiZvw3U7BEQRY1gxJUBOmhjifzNNv7pw77k+WxymnpSJNunjz+0h+C
DBUIZ3KTXJPCbkq8Gk0rioxG9zJ7Y9PQmJ1FXPUvQ2c+c58UHrL2B1vF87jjT0sR
tHF6qVrQ87dS8y04DaAEOJjIrUnFc7kRG9eq0Q6N/+XCEwn7OUASc90VnuPOfag/
dORXVGmRHBcSq1B5TXyQKHtDTMMnrplRwzkoluIJec+GoV8aGyuJTNqEnRj6UqMk
o9iB58hKWlNR+6iEYeM8lP9WAVHdcWE23/8oQiN0B046bonma1SxmdN5YbQEsRua
TLYvY4b+oNB1kjo8gbn/vaP/jXHyLo6S8qKpwSvA+VSphWlfHZL3JkSjhaIik2r0
H0DDi0Q8k3eHwSkkCFR5IPAbZ0ObKT4oSK0+U2i4p7B0aH0wF/XNIuZatvTTU2vC
zzWwCbFCMXzbaH4I5CeWnTNsVaAS1iMQRlNJUEWNOh0VI4S/gOpuFl/yHgucppVv
OYOHdqNBZJBBHyZfjYFNnZgJSuYjyBgcF+0+EDTcoLJ3ovNaHBHEn6jomzNO2k84
2oZCuP6fEpVvyIBNznstBDVGUi+bQeHbpOvh1nuWlykOxeJbQ+3F2ZXcqu/xyC/4
GWSt9p2v51kS1Tu5x1smejh6Jp6VHbqvBYTf2rsZpKRI+f1Bmx3YhrZSOosxQ3jJ
F0S24W2TjZssUiXemfrJXjGNKaGrMmuREGL2sUUoN7qwQ6GhzvEgwzm9QvNwwjh2
fLvrPVo39J77aeQdncCAaBw6/pbdhnfTXIZMrdUfuKT2ZUvL5pjlAfALcZgPpQZH
V2QDf4m/TIZVobSKGBnh7XOim4ny8iLSwVxznxsHurH/zFh9dOd4eN20E5MiDBXg
2+JC4gMrHaox6g+y3oVrB0S3K4n1yaUIbQWzCgKpxbxgmU7Nino9585ZKPitT8Fo
Qrb5v/hKm+XUh8C+HjitDmptrCHXQUxQcvbLRsYxDpl08c+Pp4C5U+SHvb/xqfmM
8dlhAyE+Lz8Zz30Xd7Tj+0BA+adkcvEy34UaOaZRHyX1eiXAT+cXuMoRaBrMiNZw
PdBBwS7OAzpW8pmRnBhJuDj+M31zmVITgQHqF6hZfIWd5JjL6Vg15oRO4uVQUQOx
6ry4XcYeM6TSU1KAQMGy7m/IEDKPxHzqWiMcyVmfC9hR3LYud/i75U1RW4bAZ1MW
KMpqnGDyB0eFKk3u8VPyiY4OIYyafbVvN+bf3UYI5VHJDco7k74gHMM/mBWPR7bI
lZPLmgWERkqa6S0JCBIQcWa4ndv6uMoRT2l4h8RTVMO31mkPqyxAVp8MYgHl98V6
Hx7JBtCZ+lro05qCbWPUITPWgKuNuoaKaT44vX1FRe4NRK7q6jrYlH25k5zfkMAt
6pi0RK4jRbSP+FL9Kyh91mmvbxh5ycsgsSlSpLhSiqfVQIuWUSEYqG2k64fxhmim
xkMlJdvcQISCcRHCVOxq8KWF0HYGB/aUZUDe8Kmq3svaC0YJE8HpXm/j17RXZOmE
mGTmH0M/a1C8q3AtXUdfRYZ8YY00AglQrrZdLZnKQG55mR7/DUz+hV0CdAk8qeDT
9WxvqvTdp/QKdjV6jPoX4TbYYlx1imUUcF0k3JMjG72Zauf0fer1to32F3cBjps0
5Iu7R5KsUlBAECSM4uFCBpzoNhgpnNgH4hEDGwXe6e4ycO57L8nDwjvzpZ83W22Q
M/+uDjecP2j21ANlpewCb3Qs0Agahzq8iRRQxihSbxaqmTA8ey8VU8OaGVpcTbZF
sB+U42M/f5HxCN0XsF4N+BAsxrr2i6kQaoxir2nOeATVb2aF+TXbm1unEonXS3Vw
rZgzr1lpcbwaOmDX8H3zXIIuhRIlcmsfb1wgFa1gFMZTHIHaGxSTTLRhcqo91NfD
PcJY3hhIDg88l1KYKu/wKPjhmevWSViDgJA3lQGtgbnfxjoAiAUFdkZc3wA9UqBl
frZG1TCk+DEskDUiRc0XtIvWybW9ayJKDJQ/qQxavMKMxaeTK3zY3F4tyjQpCvUL
6xzFzzoHmyb+NY/wmqYZ4XSSqwBXA68HSYMdYsJtmtMzUaWOH8H+7vsnNC2HDlEE
NF+uBLbq/3dhb7p8wptyH5PGQ5XN5dYE8p+/hIuADpO4RlnwGXfuC1JD4lIlxOJK
H9CrnR0eszaCw/8lQD7pf6kjnCVdlEPE3CFUBwTg5PKJbJw/Oh10g8MB+Hz2eH01
DfOMazQn+auhIwY+W/w8kRb0ikon66M3OH6t44JHF+LaQkRjxcJ1CxZcbQukdXWY
X3GzQnssYARm486AEB9bQ0tS9e2QSfXUbun9UuCy84c8YzAyjR0yE4sF3OvLOJIz
mWMb3ghYl2nYDHt6qTMCv7sjjHc8FBi8pDfOnChA+Jpq3LUXY09X2+viCh4g9zI0
tHht01GOw145XeTFoja+xIbY7Ai2x1kOcmWJASvwGcfnYOp2VYVKqtUHpPLXTqxv
QfKxQ3LpoDrneaY5YqIy5Np35qEpciP45R67MCNaHTmGTIi8TIhV2aV5BuQZMN9K
wEQ10wYLJpDfzBFvP4yhOwXWPsxV0AkH6ike3xmOYwoXbySq4mbt+wy7tw/z+J9G
udQQPSZDc+pQEr3TJM8iLjGqIbuRagD3q5YGAEkkZ+jBqBkvTykoeA+pnYIzjk/I
3jiZMxEPL3CxDNpZA4npMLK/uovOpRTQDTrehotFs/UwkFN6DFK6v0oPUax4EXcd
sX3Epox3LnQmQNXfIfjb8/w0V4Dp4QMqKxIb5PwFraiYQ9tZcaKR4kD3CIBFtmvg
4MUKAhfTP1kS/GLf+N9NRRWPZzDSNp5bFYp8m8f/z/MBMNI1PAYVupuQ8DKSQGSA
y1n16XtlPFO5JAjzwyZ9uac53zxR7AuQ4j7xt5MqDT+zWh+rC/9eKkNTGfc644tq
bjm9ICxHRerYWYcle4jIM+ycDo4Dw4qEbvvoo4gbpaCuZ+L3C7R+1Jb4u68YJYLx
HD1kf37lpiCQRQzfSAXmoMwIsGw7UdAxRWPEQkHdaDj+NGLUHDRqpa7JbC3ES9pA
980cCailerBQj1kI5Ip/Eu/4JZA1icOJI2bkB+eBzts/to16mlwTHsubo8Zyxjgy
t82GaILrEe02oL+i5L/JnPG7Na+T9w6ZWuCWHRX2d5rW/0jCxQkZSsUckZImmOyC
KIROWYgecMznOVI7o/x8CLMyKbfo87wgLvVLlzuL2goE1ArDV8lwOA0JsdSPUHab
81b1c5itawjdKXwB4iV0oV+qwBnhxpO+ANhPBBjEPgfv9+8vbw+g+LrjpA9tTrRJ
1PUT7/PEILKhDDhDFhBpUnAxd+FNGV1E0Ab1TCyOZXxoc0VT8ypxxrY2K5vrGLCJ
Zyr1FzR99QcMtBTxNrihBP/FwRcwoD6ApS3siCOUvGr4FJyXBUxyi5ah5uUWmuoS
aq+u1H2F2AsowUUl1P2T0bPdf7b57DF3Trj82yl6ARcHzeAk19B7Z3tSTs91/e9k
pEc9BhlkbIS0H1wJ8+12hYCNTgDBrkgBvsOQsplhka1Qvjs1cOGCfx8B11vSL5AG
UL63MfzTvPSDedDCog8FoJCvOiu31dVf46liuyyF3DCkHd3p4ZElPpTNhXOwcerK
Mc+bGpOEuHE5SLG58q1ieUomaNeGYLR9mBRnXWeq69Eh37eNnh3wPvrmoCqgWSuY
3wSKFMfmTHetq5kifKsPt1qjPXytk1V/pNS4K26+s1IL9gUXiVxt7ZCPgJLYiIb5
mKBdY1Xkz55qs/bXXayReR6m3pJGlSe9fUapv5EHpM83eV9NzR0HJC18z5U8NpZq
HeYajqO4BUC3EE7/8vd8/GpDFWWmHWjhR00porJH2h8sPSmGlw3UAqGmMZY1mSeX
6REA+ygh2gmtZc2q7vh2Ts7HMV/VO76HC1oU9SK+CE8bLtXcX6e+Tjt3l0rhNDNq
qi1I1pQPaTuZtjGUq+dOkU/duKxdVyvuGhiiCesjugedAU8Gy0/JQyNIPkO+48te
ofxrWLU1IXt1XJFJ3Q8/zXPnMdh5DMqSaSV/HcKgO6roJIcE9zUjvnmUctOmreTU
jQgqknbVqezfLBrcEUJnRvBseDd6mWfutY5h7F7kiV9RLIUjAmzdjmQsdp0gY/lx
XuCtEBXp/U1d+sFPgApQIf87X+02VkUxJnH+Xcc04IN6f49iXplDTrmCCGgihbeR
pv86O9HoICo1Y7lfV0uuk5mdSNGxOA/cP3II9UDI6qDF+kmGjCJVE0OjtmUskUSn
hXMNOUCJ5wRmAwIide6c7IjxaalonB2OqGYmuCayLHudFv7TktPmCjSZDosi2ZLE
7+Z2hqKr8knRhnDPPke3EF1Bq8vi4oxoLy6uWWARL2Tj/Nv5qdxt5Z1PW/O2ZO9F
VL59ZlDsdzlFdI4IBX5oBUg6KU2h3Q0/HtVSEIeM6t3uKYFTDAIsNyCY5WezE0jj
FRRrC+m7Dh+UwlBKHtEwAngV/7ses6w/hCHjBfO0poYV69pD+6O91LYIlRuSSI7u
DViIBcyAW7x2bqZyGRFNuDVUWwaflnPXmlZb6G+tRuKITGRhlRI9PV5TpVBFyyBh
F71Lg8va9wVszHolS6oVes9p+u4xRQj7SZnxguh6URUM+IPtUKHEHTZfBPxJEJOB
dBRikKOoCSnn46zjLdOi4LGk+Gh7g8bh0voek9mms89gMX9yNld4Hgr1L0idbAhJ
NztOyWSnBjXS0mLW3aHWnFAKb9YdAhhgLFE6E584iN/7oTfXUkqTQIkbe++es/7H
DOa3wgfDndvLyAg5Jd3/jlAk0zp57xrlZiFfselWUOTPt9BH7GFl+CqJXstqSQ6K
bM17n430LTUSlzZVM+AP7b8jbr8/L6Zk2lIiLK9TTWXwKG1xYvyGHZRW3AuetxI6
4sE5n9xur2Xm5tsKqwS86TNo+20DkzoQGJc98/opz/lragBHLhQPnS5Azt99MOal
T+WYQ4meqhtCF1AGNXuj1jgYAAZM77AHQPYVnG3XVTGRSih69C8j/8yuB+sqfxbh
tRfTPqSF1+YqxvHpa4moJbB8iQkqGQ3gWDJROZdACiNxDGNx6O3mTkFetybc3c3w
f5l5Gv8Hr7+UZyi2rUWBhCPAb+G8zHx5U7DIsNWp+YmzUWXnf9Jrp0cyQsoXPKHQ
Qp3BvjywHbPttnCMUbMG+3GU9R0JiOMwoIwbm2Ruy57LHtpHMJEfXfsthCagHpxP
8fa8trTWIaiNAS+tKSf/DTIBLoGyDxZQJZJTWpQuppOWGsyhQmyoinTpJeleO7og
DaBY8cGf4IHKMYKovb8VvjyNQPD0uCMJgpL6HUjU+ItMy+nkoe6gULjGrgzZxc59
gVNMCQvyHN1KRnUZULAZjL+eh2jBKAJMDp6RgAG34R4/mgLzjx3Dma82dj5kafpX
lXIfMm9tHF1F1riIT8r48nieHORx4dz2G7tT5Fh678ThiBa+43QCFwlkBdaazHOK
E6b8rHDq11co4EVG5ut6KfivyVLT7gq6iwUlA0qalGicwMc64QNLg/2Wy+lm6F4F
4BqA/8K48Pf3JU5XUYgMJl+YGPnUyi/wod8rZUe1bKPrSUINdEmAFeytHjeS0LMa
CbWICx53uorJUgFakF586Zp+zBwRB3F51TCIjY7jWaac69NIZHhVh++P+wwj6MiU
dGxfCYmbx+7JJz+Q1/sUtg3mmfcb07Z3qu1XL0URDuaJTEV0qokKtD4iAVgZv7f1
GKoKM7Hygnbp/z3VpLkZU4eab71tgB6sg5EoyojlS2wL12bKhgjOGpo8ht+A7Wyn
ocqxeKc5LkeVNLN0d6pRsDlMgIzMk1YwrgE+FU05ETfreHyPgRucXWTBODQQScZq
mpIaomMa7XchRIH+wys9G7jW8qsr9L1jgzxBO/vV/t6w7mRmCRhesnt16qrfHNCm
PY04zfH9aa0rFKx4y9IFlu73v5DYCWLfyR7J4A02KYCYUsHaR4/LvL36Pd+wO7gn
0ElzrXF9ZvVbM8pdu9Ngqotl9i+xD3DXOLQCf2EbgxBF9l2zrGVJliG3F9ZaGybJ
f/KhjIa4LsqqgnOvmzU5p4RF90AfdKQ1THnLicC38RVHRc0NXrKYfvPjl4UgI/Ug
Oyu3J7aNAJ0paI5VEcl9RwvuOuD86UspRpoVKbmj09FsbHpO5uR4K+xWXLJBJMcP
AI3Y9XIOq4Qa5n1+yQ8kTF58l1ZRheDve+em2KpUyyGbc4f/wvEDXmtHkQ8yqoJK
GIbtxnRVsvQiAgih5aPo2C81C/LvO58rBBXv9Q6a36bIU52Jrnj4zLlbnqz+56zn
BsWZmRT1oqlVBNqOP83BMe+rerOCm9rBVsOBHadSV6uJVr3CYlKjd6vzH+5TjhmT
fEXCyFtvOOUSc6/9BqZqquWBt/jhkwh3zB7t2cvDckOXp5bsFOGwobeedcpFNj1P
WdMwLdd1g7XXSt9VXrAkdSkcKM3gMxpIA8Q7GFIv+gnsQx+oebcezFDqnOvWnBYt
ILDy5zh8zwl2QqERSc2dqA3k3B32rc1XdoHFsgsjowjTH98j5kqFZl6Uz8mWYZNz
hRyetrnwWKS+ICBFVlvrstXKbLrNDmYMdvL5iCPecr5llk3BbBB/f6Nvd0KFRkjb
oKXmlp0kIkyn6tCDvP0vaftI7R7ENV/BtLeMqicPH1nC3GQQOhol+OUlA+T7A7+f
Q4dYhNYw73+G/YcPE7qn4CNToWIgO7EPGlx9yPhj+Faim2xdODmZ9AiPZ9U7oUqn
kdNbXSMD3jtjwJvL1VNwH5Kopo8pjjSpwKrUwygf8DLoX3OZsRFLihBnD0WGMKWD
khJnCJh0OQlBxOKYAl4aaAk490QlmNux0a9SEjGWBuF/3YaGWlIz6S+Uds0OtIA/
QIE189ejsmc/6zf0GO92TaZUcRcAL/rZxgORrKpRnmdQyRjUPKt4c8Nzz7GT7N6q
a78F0mtBxfqiA0a6M84zQSRGdv2e4MnVnM9nfCDw22gEs8fBFqtYDg/F4TO+FJxh
8FmFZyc2Je+mrwPNhFWoCpYQ8Kvi2KlSGB7cRwMMdIP4uu2CTYjgpYRxW/EZYsEP
kNJZWJKXrNwevoOhu3hA9wGTLQ3yPMq0+r0/DKDhlRsQBv1J2X7wXkt3vgXrwNvN
4hAP7hv/WwzxgPQQe+s+DKunwMuJOGRXUNJyN4ilyTxQvFcmN+zXNNV1cOnUm3s1
hL0TY0KtkQ8JI3wOxtrXVytCuo/OAcTEM2oIKtdYZKAUjL6moPxeqs0LXp9zRx8b
qxMDsAhlvC18BwAZICt+cswB0R0Q1ee3+S8MO/5JHZClywfumdhKtPBulON834Mm
UY2EB66WSaIZz883phvw9Wt36VyPMki2eP6xuoqVFCYNtlc7gqjKZROACkzHT1sM
ii7Hl+tK0yQ48TK5ednbnL1ThPC8MlH7Iezeod6+Q8r7DLF5Uc9OUS/Lt7uokHOE
3i6GjsJX0/cNKDViukmuZoM7EW6sVsWKe9OJPyRthu/xdMUeL0Cy9/lRfApiClPW
pf+FLJjWcWE0C0/K53MOlBnMD5sN4ZyHwddnovshQH5jwWJ4B+OioSpzIBev2pmA
3IzM6lyxuOx2Gxd1k1E+BIP3UL4rwXldFexsmCRE1+dtJzuklVqNzpEv1q3MvAiX
iWMEMFz+AD2afOfrLtqpXYNiZpfZGZguNqXyxwQZxxRRzBsmZr9PwBAfYhe2o760
IDEBP3EHooudhPGqN5mlVavn/qLTrVj0ldj7zrn7zddbwSJDv9ACK1a7dEe9s5Tk
BKBx1m+y4Y94vvgxbleFv5KTELj+6c0Hz2uphVVG9Hra5TUcnSbqG8s6Zax+gQM0
POXyQ3vjnenAfTqIdvN+VRMZ5kr0xCq/KdN9o8MiFc4G9FscuGFk1+2P39MSJTCs
TSAJtQw4C6cX0RAOAOk0JWoaY6vL07Eq8S1qWfyciHzTjSb/g4Wo6nc+WVYSQF50
/KjhBpE+jwA74G/Bn/1gqUHGzpThZBK53aEe0oDuMfhPOXqbyieD6rdCmk0ETDyx
hKGsz20sL1KCCvddMDzhTrQOQ2ZRSqhPmidvQXwBjvsJ3JFEh85n/h6qhujVwd28
HU7jAMwYq5VQOEg9RsvtRP2canUr0f4QOESlRi66fkvDMEQJcESBaqbupfZUFh8v
J1TP+vzie9smUENZyeJ0TXqRaJ/D7s4rk1IWfu2x3ZrhxWmWEdneLuUlcqupYw5i
bnALzrv1om6lGVo+E7lBZImd9roM0KbSd5AZingCA3rP72r+DTKFWZT//GYsyK5R
6x2/91dcIknSoOPB/YCW29xomr1//mpVY4VSSIYjmlQjKg9Bk897Ok7pFgsNokha
dJInVKdblxzsoR9x1VzWW8o99HiNW/NmCDPJu6oCd/FkLlV6URp26/cTZz4xjYif
eSl0VyKxWb1Se55xxE3mlAAtuOEuBkf/wl97YWeUARoZjmHadxZrmfufi+lAPcmK
rfuAlfbqyGZ5NOnJWTScvUSK+anAmNBkR/wj1bFtL1j3ieNZUZThy2p0jHpS62aZ
kaY+RRzIPIf+aGDc0IU0R8tlhuj9+nQ7HdJwtShfdTGCzX9WJpi9r61lBD3dwooP
E8Wb8Kr+Uc+tgYgYK3WE00GWSgpnM6TAkk8Tjo0HH4VeuZcHNDo9HxuJ+srgdezh
rM6d2jwUAzG/cVkIaAvjojjoNAVd2NVfOlN530ChoDSeUozw3u/pAf1WYbhyjsOM
uUbe8b7kl8uOnwqGMn51kHUNTs4mIAsxsXOHhPGfXzGVNiX1hXmoVKQiWpjdj+bb
rcPV29Gpvzo28z9lidu9miL6PiGdcsv7vtKYRF34Z9fIzM4n878ksbJGgfB1tjkF
Ov6z7rEqUUnaTp4ZruYZiWCnMX9oA4BM1+l0nl7XWeA2fgdKvfWAXX76tejudxVl
jzjIoHd7UmtzhlfIEZkRhks+aBX4nsmMknmbnQ3/awdx8XPr25N7wQmIGAekGorC
X8kmqHuQuNbHOKA0l+vhIDIHShPPuMDsfrnZxwb5gV4ZtB7jYIUZJZxBzdAgSIz0
y4syx9qdQ7PA+WNv55z5VIF9KwwwIIg+nQDlBIOTLniaMt00Cz67epslHsWrO9V/
UMZgp1wKlOb8ADUIXYRnNsOzPsoKvjSu4KYO9+ssdLOhp35AHNfmQP92Gkqvwb9h
nQuzF97IN8/dPFlBZ7kOMm68KmffkH1H+VlVaIdRvbFVC1PuSnPDlCAb5xvPuF9F
6CTdoQHzl76V2sfPfs9x29C84gfOv6JQ1Cjagps3vzRdae2w6RRD3yR198Sh4iyK
7jFS9mt71sJ8bVpfpvw+9y6dqVtDBmV7eg06OpykOhmEdpoP0rv5ycTnW1ALW9NZ
OoIoYMA7r1ihHex8vWq0ewuR01oxt862Mq/o5+YhRx5x4IyJEl/qRmE2fMKT2Is9
fp4QQMn9rjA7vYSX4Iy+A+WdKsAmf4x4fdnH2yUa03cFeDFr6D2G3U9IlFkSBjh5
LVQAPj2f+cENF4RzIyWxoUft8/VGBYBhabvlD3pvdvWJVI5AHE3o3uTQQB6gQd6r
tIjMl9TXao+4bJsxjzDS9Iqb2CpuRpW/4G1ZArPV4GByNYl1fL5KNfrcX9aLAzd6
2RtUOcjNqiZSJOwoPRW6pCgNhqZd2IOhCw8IlwZEFOYAJF/dL0jb8DPJgxFslMOd
WTCZiPNlq3PCIdZUEziBX2ijlNf0Bl8NG/TxYdV2mVBPrctPECbwMXO973BhkULk
27yfFBXbPwtb1lgSMbwGOG9kIvVya8y1J3mIcw/539/Z1pNy5thcFBeJ/PNGpank
pzNZUjgOB7A3cTAHwNBxXyan9qsQi1Bv2w0/s1nYdKlIxWI+0FG4Hh4tdWYA7olk
1v9/GZSuSwjL0Cfq4yP5ki+wfy1zRfpxTTWCYA5BdI/6uoYFUMrAPEgTmOPoMbxZ
lT87fZH6PQU6WkDs5bhsGobgsnDj+QLjYwA+Szs0x2JzDbqZtxQRoq5OwZMx7S1R
b2AJMjX16JwuDLDjiaA3MVcA50YCqbHcBCPZtPrCq9kkMY9zFNQ5ledI2x7VnBWD
SIwQEkc7rC1kHI9XItl/NwHkZozZWscCeVTWeip69P5a/LS8DK2xgpbTTcTN0J1J
8XjWfj7CAb5xnd9Rx4kL5xvwC0aIUVv4koMXBspWj5UTwYz7Tfm5fMBmqkgsKxI1
NUZD8HnUeozwLQONcXvVktdUkEdjaUExni3iNqM/CDnHcqiMQQlstraSPKbRrJob
Q48eOaUDo7Sxo6o7AfXjQ2LGKnj7SGv6PwlRKJxn53gEVPgmjYHPHS8vzLvXX5+C
KZB90911S9zob7IUkfIE/StnjHMVwlFkVWl4fnXtLeIbfRHRJA6ocqA+Eu06PDxT
b5xzw4nQ+6D3i1bqnSFdbDZGBOd+FsoOLxQ4s7NVT9Bm14uJmHNT5n9uRBsMRlvD
7Gm+vDWlD38hTgc4qWfk/HYymNXCVFoLJ/p+fyU/ROt3Vm6AUrv0VclO4iopu5Xg
Z0c6WelzPrV8D+zb4z12iiakH6ryaz0TSeKrvEwy19mB+XnLaJ4HlQYe0AUQPcpx
5SgARuSTvaV1jkmniGDOsD20yfZhmD5V4jDHD0Pcg5wGVZeYS2Gj2Oam0Row9HJM
wNeGqctmQ8qJIDnZ3XMd9RyUNEaUrQ5+2ULn41FLb9/I/RgUZTCmNEj+TfKIZyNy
MJnGUBJMOO2lmylg4WqaYmp94ilVekcCABA/XpuYbeTQREppA5z7aOuJK9xC1Qge
HrDrU6TBkyckEfD6mfHy2MD+TkJzpaw7CXZMjdwOd0Oo48QR2Pq9EacYnRCVCcOj
F0bqXEDl7CuIhW1u2lahtDugnHVRi1Tp6BbNWVzax6P0scjbaoLq9eGRaP+/Az5o
AxJ2TGXWssNu/FU6IquM4ONepfAv+86uzR8w3ODgncQRq6+4daQXEGaajxOELWij
Yz4pho/vq6YWHKsmwxies35yeGs7V0xgmqfM/5S20cQA+4Cl4mrEAnuqoKAormcj
Hf276F5XBhHbMzEtDKVQ4O9nRJ37Dv4D3WFCxJPBN87gMn1oyZb4JPBHue26EeCY
PLaFA0CWFmNxpJ0i3E83Pgdisbm/FnHT9/DC1TD6VAt9zLBGhx3qUce5/hbGmYZd
pk0W2Dy3ACXqWflth+DQo7pVzxg3oo3ThhJYpvvbK3efXQow1kHwachzT53hMqzT
o502p2Q3uRAo8fJ6QBq+xTbCiT6EPSyav+TGr3gflIGqXP1+W+tKXSFfApkho4WY
nN15XdDYTo4Txxv55V0vFoFB1tN4/hHNbxuAp17KPJPVkV5PsXAFky7eXq17H/id
Qhk3uP1BvhtFp9esBNjHRTe4jLh/VTOvuPPqPVkwDhkGvN2M6WKkkiwHXuvez1c8
/R/LxasO9yBbhyeslQN2QWg6srCgSOdXsfRPDcM2CPbLcJOwYfPgbgQrYLYd4d99
gigzNnATnBLRCKMt2bfj+EirpsjtjVIBu6Hxli2dxrtlUThTSahXND3V4RHBWg0S
VlfZMsEprajDNMBCtfXDZZuUgW/Y3l1WrQC+ew8EPkC3AdnC8CbkjgreekDZUWwN
0Rfc1IRmIms9IuP9iTJNpBDRtJ0RMxd8ca4rJKqhNr6zg2k4PiVRLKxiwcfDvupl
pxo6siK3Dr3jvu5GfZ0WYmm/Us3ILd1mIxazTYYFtg2iyyk4pkgf+dVstq/dOEBW
DEH6IUJTHoRhpFcTO1b4Y9r7GfOdD4ayzH/cAGACAEBJ+bKxMduO++BdXB7jqAGL
RWj3GvrvIpgRpL0G8pe+6bEAJ4c3mscQmz0s6V3s6tfsH4e/eHOJd437mtYhH/xi
X+cys6r8LO+IsoGZX3F+6V4E7USSb8G27+osIreGC+3hAGQ87Ag+/Cbk3iYYCwCF
v05YBdXxKvMNMOnpf1Sf51bzn1lrOESj+Decd3SOuaCQbzRvVXdJXK3+uyeeMb+T
VDzoJgiAmE4tPPEiLcOVXwsG1tIiC4QOYEo2veyUeu7rnSOVZa0h47L6Oohtur99
KSl3SQ+S4bEIZ9scYNRMRG0RtlN3Rvn18w4skMiFQVfVAoi13mHGa0e+PW/sDgpN
S8jzjmeeN8wL7tBXkGy0e8EvxguF4lVwnQHDASlfysrnEvnOsyIgJuVgbF7Db6q6
IiHE88/1skJYpXpwBxl0E+VJGC2xz9lkFpIjfUB9ojXP7oXlJU/zxGMTnEBckPq7
JkxtKkjlFSzhV4MkUhLlvxKDU0LQ+kiA4YcN5ZbrisSlYuFGnMuDqKLRo+OtR/37
xRLiKRxAbDqP8FfWifKSucp+PA4D3hMkGbBjdT8vsAVOOKh+OYLm5JUDod0YZfRF
4z7RMcNV8yyYE5m8v7QhSWYQWRLNZkMrQz6cYqE9q9zWWYngMa7fSbxEgK9EfoBm
1iBSQOD32WsqNI5pjis2OG2ezn9wP28yTGPHSUxCyDjAPs94USLKECM6R7WU5Ov5
m3jwxwaiKUXt8CmXRE+4wb6pgCy1RpRAqorn2BJFHLS+HkiWQrEv/tpuZYH1ohUy
AtaI8njBnCPqiytVX48dtQ5NszRzUK8WgWG5QRhTVp76mAUaV/nBAOLF0HRg5z8f
8dWP7MY+sUFKMoShXv7Vz/P5KC1+zGttd2XgFXxprsyjoOlaPi2iU/o5tUY09LFx
+8YCczKZT/qECk/oUWaIAZxPvHU1rHltFRcMHw2f3EDq2EkO9qFNh0qZIvTdXSmY
3XJNxMmfsTIhgsYKy9kGRPNGC6L9lyVtK82OvIUqIj4zpju88a0WIjk8zEsr8OzH
/rDG9MmPwZNrOxeBGletEgFIleF9D+/g0vc9f3q54DnrPJ1hD7rUsU4oWyBdowpI
rVaYjCKmOuGlbA945fWDWtOfjy7l/p9sxgFyV5Q05B3RA8wi9zpIzntdsYDHEZAM
lSdQNLtizzYlwuve1nU/G2uDzzbTu2UESu6+kf8VbhBBsKv5dbHHUTy1yKS7vBIj
CmxiqaoWGEeirMO6AeGFq9wheTHEmIreN/Wlty5lTwFakFKRPf8/cpvlcVbLdyTW
IFSVDWF43oDcN16wnAyeU5U+NzgLGqaT/qvxk6G4TLL/2tL05boxX+sYWuu7yyz2
azEB0C1ASZIfQNPzBjuCHd8/M9uyrEDEhTFf7po6nGsZlSR9dnpQJ8Cogoh8dElA
BH9dTHuaEOmJTCKVIPNfWA0fFp+ZIDAsQehEiJ6Ab1FRVGYpHGohsQyblOIxn0i1
E1e4UfUI6D309FCYWATKYJfjCOzWmlWZbQITKjmSXjhTSIABPrgHxyoFAEA/2Y+2
Out91MoeUMymWZzhiXpKLK8+lKH351GUTn9vGEyuPHGsFQlDz6nhjh67Z7rgAl+b
oJYltB3RE0VRjvRfKyU/JM975TfkIg6tCT7FAyPbb4VaXUOkGxnGkYBn8+DsWH5z
aCFtnr3pu+2AVyYoHDvKrbpNXvSONpAfewwA0dG2BQJlzHvg7AxxID1PfMNWv2ny
PCpIO29EIocBixHyKefgRsfaCUKnXRcx/uMUJb8jSIwLpa3ktRYvMVz1XQPMHYPt
OyxCbbJN0EWw3d9fQmh2LoXu2fJNHIq3yak0GpVYG94b26hSJ2p+AFDI7itTyTxT
8llgVN/OXuLAWDSRuyu48k4HOYwcalY3md4jgkdsNmcPoGa5hlLe6fWwWan6z8Za
NHuL8RuyJlnJF/H7XxJ3i4UMhJ8ILuusoavT2/LVbtNY76S25HUAp2Kv33QFNKw+
MEwqVbvgrs4zMiqFngYc5924riOt2fcjqyhHQ8XPGGymX7GwCKZMkC9Mihx6mujj
AVTuy9DIl/nsjQhh6GiIS/36HJxn/HH+BqJ1l7KFM7rEdlhSDFqQiFZeBABaj+x4
ILtFqpBK+x9Q09pATqb/bZGQJGB5JW8/qhpHDyiarvO+nITvj6pIIwdBnSL89e22
BL2S0K1YuHnt3MDRb1efNAEwWH6iNQAN6TNFG+hPIWQJy/ZeWXSmaIBbotFFK1Gx
FUFGVQRuV4Trzv7zCWsM+b+00YjI2RsAYnsKiMa+WctaKPf3GGW6UHSSIe8ZsSH2
9ipCrtjA/rfN3tSZ7dgKVIn/G4DFm5JJ17vKGxy8qyRceNg1MFmxgtYxqgRLaMYZ
RhFjRlLUW97JcDKCY3rYIwGUNlXbWDUGlcfBE3Q3zRx/1QR0fxbCO/YlmpgVYPZ5
wAqlMdNEQU3OEU4Bvf4aTWsf2sa8hg6cYVXaQDFbShvAsMSZ4bNErcSwBS5mQz0+
I8K8o/WMOb4mTpnatLzPKWZeAMgJFX6E/jsUeF5Hf/S0z6RXtVj7AnEuSJo6ew/9
g/m1kpi+S6vhBmu3HDm7ltUTYLpE9/4ibDcSvXKwl/3eanxX/tv+gLBd1pSNMnE2
EdC/0VRwGqAuuRV8dGXgJ428mCRvudqgIaukmtL1P7QiRfqFq/2xnwHqX8hheRtp
RkO+YQiUpOM0ChOjeJvvKkgG5m5iezvyQ68BrTHKSiIEsC2h5wNfUtD9Y5OCK7ca
Re5mi38zEJSA4h3/quT96LXfeX+YxzInP/X6mf+n8aDKxl0IbZbc0O1f6QAMURm5
rKsOVBaEDOhRY4KgcJVr39fxeVnzOaVeid39on/UqlcGrJygBREmIEewSHrHg2AB
xv/txV+NVFAmM9zFHtVRLmNKr/svlDReQtKCVV50WxiMZvKiTPv7mjMk8QgBEtOT
hSeEeuxtHQkEMzX0nU2Q3xOWG/RLEQKByP3iKjfghl+mKByyNvR0/ugCOH3psxPN
92eVNd4erVfY2lhFkwOhb8vovRz3tHlyPooZ7/D32rLYFvjs2KSCixLNykb3Kyu3
VEZr5KHYqmH1zoSWTSI/MjD89yqDxuGGcxm1AgeH0W7Mj6KQDvLuyb8GlGoDv5o0
aZOUfQ1Gs7nD4hh4esbBJ65TilEEYGLLnkhTmpO6liNMLqdS6/OLKQkQHVEfRUP+
FED4vHOT0nq9MFBAS7dDaCEe9zQH4gtaHOFWvpUqxViQOLx+xCzcli3cjrhd/NUj
PNnfSEH7siW4bR2kaMvCwBlhXKe9n6QeA1rJNAj6PLvAsgjZmKStTiAFMNyARZez
00P1iL6+d6crajCQFBseYTfwxVahm1ZAnfiZNZwavMoRKBbAVW6p6RH6KAmjYw2e
WMVa+f7gj1SSxNKZSwbvs+edRW/3GbY+f1JMn5BpDJMfp64xzTkQrXVPa3E7sL9o
CNPvvq9ndpWqF1pB1ZeyCEDijwB4t4mDEtdb+pXjcJo6j1H2K7rKKtLL59OGv+Ud
pfsghnGWug78nKEyIWLOizxDC+OYVCscXUnIy0VeBi9jUi5FQSqu+1cXqS4SZ32h
yA5VBmOhUBUotkAxd1XaQW3hAZQPEf+mxzSqganA8YgIL/ayzB1Fstqsd71Ujgtd
eQCT3LCj8XVvPDk66sO8Zh7kx1LHdpY6w1rdA4A8ka/CiF4bFj4p6LvTHLQhNgsv
Axz8s+SwcQBkdtuo1SU9AQg/J3Tu/gZzLmF+z1SQK5kDPHGMiBYbX2twQsBZeVxC
XocVj1kySSaQZT3Jb3F1qwZamO4UOwkIEosRSOvT4d7u5xDO6YKbLJPxab2ZWIBo
fvu9XRTOAEfpROyJEHMajT3BkKedwsUkuVdNZzW+Y6ZAELnzyOh48C2pGEAu0ay8
nuLxzgLrQbPOkN4mTskdahYylc9wsGZfshJJM3+wUsIusRnF02dHZ74WLMIk/e0x
n9/wSlaH0QU/oo8ye464D8P7cq2x90Ndci7WbkqvfxLO4PeiGwYvH/Qcm2Lz96CY
DUvV+oi23aCgE4l4QkJ+PLCibZMRV8qH0MEL6ftFQYXXyxs/i2kiuez1iH9M/PHr
oYWE10csz2HM/4AaeLSKLPjqGYDtzdUN4w4z91ofb33z280ttvtnP6CcqrwXnQad
y7i6Rw6HElE4QSoYO54i8wi3MuXM2uY0VqPoTRfOLDahoipEPuw5+uHz5to1fGkf
7Vov61wsmRp7XsrxJ19SqYO5N92DOSQXD3m4FluRismk/o8lWyXmPnZF/UQTl5sV
PsYrIGPl2A4VUUkEykrjFxvwk+Ck2faSWBPmcSYs+w0fLwz+s3zIy5FBC0sbR5BO
gojj8j4dVrP1W2//RBAkGE7NwQ9NqizID5lTt7ar6Xn0TwZARb8fybDpephRgV7O
EyYyB1e5e/vACKngIBggBWx2Aivi3mEpHIM+ui5IxwkQ+9FfNzWYSo7zzXR6PBBA
SP1l3Fj9NymbzysuwTQxQWXPUh19PH1WuCiKBjnPAbZoPrC5NgZ23xNOx3qaHXLq
GPDZfCVWNWeEbfbv5CAwTvS++S9i38DF1AJSzBxYDDQm6EyfOljj1fNKuy7NFkcT
Md9wxtCPthgKuN7NpZXXisJHc2esmX/GcTn8J2TNtfAUt0lRB8Fbd4p+GKGpRuXF
Kf1i/lVG1M7gOpoKOLkoKmWlmaSeCRSd7N+nFGi/LOosYdWN3Of1lxivsQWcG04J
FY1hTEMMg++KOJosWDL3e+z2a/h7jRVcWe3Brqw+k+ti4FtZL3vl+NM+/nnLfwuC
zE6CSvaot6WOxZzkYAevCHdNITXSSlq/vigc9uHjAUgUlFnGOU1nNKvRZ0deTSqM
ymsg35jLd1BtdWrBdWUqWreD4YbnDgSFfVfVqMKWac2X7KsCvzCwgPeiPkL6Fg4/
LN4wDeQu81N8FpJWY+JTHELaqdkt4X1ttq/7qeClX8jD2Ia+gUb7gNssdAf4lSdd
S8OI06gIBl+zmpie3BJmT91NRouw1x7CBVG6vOcVkhDoQ70UhKF52PnU1s7N4NaG
U+WaBZ2ED2MPRSvrYFBfeGSSjcZUvPejAQYUEmTAQGp8hdSr67jie0TD8dJIu+hv
j9rJ9/F/gC1ksaO08Gkma8vJEPjFy/5AQcg6j9tLGVy1Y+oE4t6Om3TQv0nq45Fg
75oYDtQ7SFAXLPoDGGmcDz9c/wz6v/xvuAQOQ7WZMJLtD3uU/A6ckCJkv0m/Q7/P
hb5ybF3DGV+7foVWec/6PijEe98QNOqYyTHCSuAF720d3TDln5mbG7AoiWKlhi/l
LQwD68c6onByAkVeColvIOKWZP7AxcK7eKaXwhbDDK/CX9pjg5uBzvG9JNJyqgnx
JkTxf/VwUke0oXorSrtVxQNwbD22Gu+PVBQjwmF6gwud1g6wKV91ss6HJ++uTgPI
Pbo8QMVNUV41qCQBhEyfGZV8ncpixOSdpL1gvvhKWYVaqqvBFWdeMODUMWP1uIUx
BuU1c+w6ccmQvkSWvb5ri3In3PsFa7cjGW8DotMkDIkqw4GwXBPurinRYNnh5Yqn
aSelbmoLoDizdBunEhj6oollGssT9hgHNUx98Qf5v9z/hStoh+0lZ9Y0nMMImdn2
0LDkfeS2E8lDgylVnTYHmpi7hK47dXURzkgAXhaTXjQoXRfFqNIBZMmb9yLT20b0
Pukpd6kqQCTU04kVWPso36Rbe0spRgp5NX0qA4O22SBQJK//AVSjWMekDee2sDrk
s7PAM2X6nVxdTQzwevZ0tDfZigaqmU9JyxpTVrbZKW1qAFfmqaVyFV0iqVpxet/2
EX/vzadtGR34rxV4J+A614MDyWQRmBdlIxn0igddFFWe89E2t7ClUdcJ/1QziiRL
Gfv8sohGYYR9UScmiXvXHhBd9rHymbyc9psZrhrOmvf+A2EfgeF1D31bt22ceTpY
CqajGOZvCQadzgr1OZISsglcQjU24WCCgtVgY6iIQZxeeGvMPdn1Hhmjm8Szkn4n
nMu144BmD8aUIdoenj3lWL3eC/qqzntXikH2jDdNyW+or8E6qNYcNYAQk6X9P5yV
HPVvAlkGr3l2CPTQpwRA0RIPesqKvWg62VcLxUjNyg5nMVvOYxKw8lhmD9Kxvala
96zY5KsJ5UFUxVkbgWMkxsWR74yx9kgiiHrxboDZfI/4P3Tc5wISfssQ0GJZH0Qm
jnkHnWsuSbLLeOA0qwSMMNNEHXw19WGi+H5fEThM5Wpl6/BOibrGvYwahpek9oHR
hjNcF0JI7FBhzT66x5WJMzt+9KYScOK8yPMcfVB5phomDPZSoQNITxKMmIV1DrN2
nuOEuBA9byrCnlTTKu3N+RdzskNC/bWA5taGBZJJaQ2OrkZc7/HgAtlJKA1CubHd
+afBM2oHhPBGl0s98jjDD3O/WEqdPo8OivSTNf+s/R/v5rl1l2BkxCqGxL5xBBQT
4BA+yBNKWBgRJ1yz8lE40a2ubPwtPImmmMFlvf0hjFMG9K5FHOWdFRC8nDfpFb4g
6mPoDzTOxVOvJ2jqdOa9I0tqCq0kBW2xDsqzF87ht/KHdnHgy6rc3GjO30dsNpeB
YZmT6lhFMYUjL9VC0qQcpHxGQNt/kk1y/AHHHjB/Pxx8P8HbbpFrqO4lAlNTa0WQ
rVzTAMoF9MMx7cKr3i44c8BZkcJa6cfkLgGVS5OYE/BG1NJS3a7AzW3082IAoPN1
a1OzSUQVBbt0DVdEs6xMbHhCjWxH7pA7KNzK9NbVxtsqhWxri+xwn/VtmMBOGmpM
A7Sy3AJ9bb06MMYGmFGW/9M6OZC0DksUqo5+LSX370YdgmkFsJQAr2xGxTFWgkNh
fhvfz+ECZioeeqxY+xNtOEsHSkOQ+1GrsX4zsbgRR6CUGN47Oagtkpcfe3sS3fSS
Uy4s4K84IVmQxOMv9qwSDxT6YIjjd7jyyzpquDHHMb9OgToZBOIulo67FQaFJsFp
DH4Q+dW+vXZiMSrIR1OzXTDx2StnDKjpw4Gn1yFiZBR2MD0S/9UGLJ3r0XUBbzrv
SY4m017x0vwjTSVBY2QPJujEoAsMegCyO9w9c4RyDZMEBtIB5lJzBVwiXuTfIUex
binedprALhPQcmMC3brjORqaWUQFP+ibC+x/vtVqU7iDT7TsNQ62gZCDYPKPByEt
nfQDn50x5PIE3kXJl/OiTvY5qH2smJNEdaH6+/sit1hd1ALAqOHO81yBX4toOlbi
tn8jZl3sV6twbMfEg1GTbiCv31AKHOsa+BKlKctG5CoLLVd/zsvLNk+wQvAdVpMR
fyOnuXapOj9YTrvgCNgV/DyHXKsF5Vv7Kusz12MbS1fgy8/RMDyzeU6npgD1Dn+y
xvP5w2LkzdKZwR80nRSEAuxwC/imIpGzIA+7cw3PKszRYSSAXQAPbfg1vpXZYizd
1Yx9Z/ilhYd3u/N3z5G2GJDy5nLjoa7Wo49f4OTGuw6qm8m69bjncQTGzxWbggq9
2by8WxsvRmspz8JqvFwg5myCyWZu1/EJ71zR96ltv1lT3tLbTPWSvh7gB7UhBpu9
rJXx0dUuca5uDkKO5kSA3MznkfgQo+QwYekXnd+rLqw1JSd89eqwCoXS7H1he4hn
UWArm4u63nKi1ryLvba72IbDNpb8HQPRl9amugJh7ymcClmEYFoiXUFbDtQov4Z8
y2/xVmweZ0EpY1N/nA+xWGg7/PmtNfxjn7cvMNFAQ2xXz3WvaAS7wUZ6v5f6gkCf
kuRyaTtfiwXbj0M01G6OX0ZeqARjmvRQSWJQPW74M+32xx8pOLQLa8ywLA+V2ICR
wCnlLMGNubazDJHVtWY25Nwp0LECRGVLnk6+eP2JoQ0NDgCL1tcZYbnMloDljDlo
Ny4sDQ5SFjY5qOClFq9D/DfiEp576pfZNOxkMpAHuK84kQgInV6bK5ue3CWbJWqC
D3fEhuayoO4JjMriKZHJPmy3A72bbUC8MDm59/Qyls+fqCEPuf0OoFRT82V3pRf+
aCWGFcnbH17cmVELk5YplnSRH0Uh3Pfem6Cwo8sAgDGNNfJRR2cogpg1SpJoxVva
aXlC89BfZ8nwuFtFYj6G1vafRDyEsB0ptQe2Wk2w9LEjxg2DSTUB19TCP3qhNQrd
pNAPQ4lXnbajxMQo7/4iRf84f5Laq9IPiE3vDl8qhJvktQm6Tva0LpMdfNZqVey+
Z/St4Xc3N2HJfjEWZohgCh7sdPNM9eE4pxVQU8oHgpiUUFTd/LkmuVxbXfqiMe2x
gB/X4CISHeLu8whVUBJ5KLv0nDO22P+mMx9WR9F9bCQ6Th9yhWrnuRg/WEm1GnrD
fPn2jnLCx8xHKJcnnaAVv507leBj0r/UrgtECjO0KG9IDaWMWLiKDpnjpt/Z1jDz
Jt7FUIOmS45EmgYSJTg7nSchye0FqcBvh6enAqX1fYvwDb3viS9JW8APZ73j7Vwa
ew43H7+0IkT4P/LaLkfJkN2xzZSNQwMlIuYrRlYOZRa4W1dcUYYoo0V5gms8V5rT
qgmOGNu8BNxMVcehuk4aKR5C0cdimc10w/iY9SRZKkTRem0LZebsGPQNCx+bYfWe
y16KETgN8klBSibuImFYMZ66kHDfV39N+BlSM7aHlyM1XVumnXTfL/7BLODc+Ggw
17ehT7MhFSlKEcviNMB3deXYPPPrHKf2pqSpqBxxwiFsIyV8vwCFVXhbm12umxwa
suf9ANEegXdOpzt9euAKSkG1TuUR2f4CnW8tVjsOfDo8B/Vl7v5f3PASlLXXHhYF
N6DJQQVMTjgijfDlBgAZG30znHN1Qj7qTTAkoRHI+v9nmnAyeldXKpDr78Gd6+z6
DQFIKYQE16FoGQz1cRpDUBMY1YJokEWHeQ8m3FWb2ydFKAaO4wsDxcULBS4NA8xa
nfmTnI49yK6eu6yoUB7c/LcZWDaxrHY9llhbl7AAj3VnvzYXKAi9hfkqHMW3SG+o
ZnG4BvvGGfr20LjL5OzMl3wt7gMR9gs0j5FCaGlBgRIq+pzpET0f+9vFfjsjpKlM
iw8CGC4WhxGOiSB9trZ7SQh50fCif8co75FXg5E/3NuKR2dz5KaMvDjdlsjT1hmV
RUe13iBe3jm+5fiXoixFlutXfag4BLj4jzmLfL1l0rtU2PMy/124XZ9VTNLS6rg/
9+w/4H3HFcqSVxHG3MfC5XZ6wUcYoZAcwX/ORjfo8oKEr4rVKnH7Q7/xFlb8miab
llN3LcxiXM1xtlAOw8bBPJ+SIge30rMiVHX1lLQb7IJryfCyZdBo4k3PDZiNBfNa
H9V5+LjvwvEo/0qW63atzW0sAr2Cw70yhY5xEk0Am/7Y7AXCrHrGmf62+61F+zBM
tQb4CSlt1yZH+3EmGFo1M6mVAsgFIBRcCEobnnLHTg9Qab7s0MrlCSD/SOLqjNIp
KdlAH4RNLkZdeuQkE59/xSc1IMZei+KL99axwa0/V/h/EuIkxhcApf5erw39bxnB
rT0uxfNnz1/EOnO4FJHvV4TTT/5LXDWHS6JitnKWWU+6njMpVToa5Ga3AVKSdIdb
ixcyukpLB3ad/P+2MqG19DlLDJg7fyG+LLLVYE203qWzErDbANjDwCddoa1yYLyP
nKlu69M4g51upilj5VO37l61XC/O0KDHgyHBFRoSoZYZuaiy5p43ejFZMkWyIFsU
fdmZ5ST15As3rqOLgKCFdOME/UWcf/lWclFswpJW0pbta+EQVkNMlCRHhnIeAe9M
DMIdB1NWSK0eShMl5theuwkSthiXbZhnJ/dXlsDzxpi7PLEKwUD4V/cDMxQ/Csce
zF+JmKR950y7bgkVRUdfH0Zimy6RmFaS6bReHrXUebf39+IT62G6pD3Wm9eftUed
rHEHnwZWC4+TXpkNLMLPAHtULg5JuG/nJhKZJ4r+m8LRDEdWTOGHBvWiUdmrRdzy
sugzF4PfRvsy0Xwv+vOG6cl1LEJBXAqqNaS0k8rr8CuIFEXM4YvShXB1WwYmTRHN
SvdIQ/E00VSuQFSD0JHQz4mHKYkVeUNQx5OOZ+9uxaplDE0R/wItuG9TrQ+cZiS/
cqEKRxvzW8ucGXYHFM+qEfS0TXiC7vp42Ujy7HvrsnGYzOd8jA72CUqPCNPQvlLe
gyyJhz2hIlSLQDOnjjnqrMRKZRgDFsytUrxezTz8CZ6Txopqwp8NmhFCmwdsCwTw
1llsdIAyZJzgtpJM6+xmrw++EjdzIDKCYUbFO41XR1SvbxIQt9r2jxgzGsENIpQz
lMMiZi7uBoWGjSgLdM8ddv73QwNdNOKhT2VTN/mSimbw46WhtnyiwccMc7MyVY2+
LeBjyZNoQ0BZne4SDh6289N8siNrkCmW/wYcPjUomh1EjAvX0I2igkpvSao0WOPZ
xM2SunfmgV0aL1PEzmIOOEEuQNMWoJVrhjOyQzoP5df9IpqgsGjl6zD+cdUaxDEK
OlcFzfkjFxy0er/7ZPSphx/6Q5G4OedY7WZkU4N4pammII9ULWFgvuF5EeHf2AXE
K/I1HWrObO8g/pdiZ1+iIVjD0egVZGJwXVOycyPHIyrZJoq2CvtNmXGJeSanb8rE
S+Dl+cWcRtFXpY5o1fwtU2NtS/qecXiOJQZ+4YSKySZ7uQXHK5W/N24x4jRZFNb0
m5AVLnoQGJdaVb/vdgepdok1yN6Z8ODCngKAEmKgsd6Prh8k8ccEa62WZ/7NMEfL
QqZJpjTEeKBXeqmZ0VCL1+ekT2fImv/67dyjUGq02ssGtiM21BDWF8EIw4Rl/b99
aVobTIfLmlN1HTJ2ExOiSw5FLCqM9E8RT5vmnHsnIVivzhldEdTAgt1lOgoiqa5k
v8UbNbgTp5IoZ9DOCicY6JBlctsXL1YEygDgIBWH+2797r8WnnkO2pbq8CQNsPTi
U/RH9D9r3Ffht/GLmFQrnTHLu2wbxUa7NBD4qkmR8J2wtK93kdNreXYn//nrHQ2A
bynv19iBKKYLV9tzTgxlSzqysyT79qwOsoe4MwNFXHNup90AyzIYdOHtZOyAHnMQ
/U5eW5Ppq7QjsL3YOXnwc9ypPcPLNynNsoo2rucewtO1jH+sPco8JkqpsjSUFLr7
BLfG96S41grVW7039e3xJJx92bYDuUI37aJakxX+lFGCDSPGH3Y3tuqGQtzSHG6u
Wkib1Z9e0iyy5ycI77G4/cMuj2FHB7yGURJem/xldpHDc+HAtmuhoQBvYZzdFew8
AcsmLoDvqEmqkYCzdLOFbwfDYnuhjMZzrweKKMXYbjoIyaVJlks0hKPdRCsnTt61
v5Qeooz6X778G3KLu+gE/jwbMqzbimu3NufL3VuMRQXy3qI5vb3t33OyD3FXH1di
Bjda4wQ/iulFk6KEY3cMHeRMrVDSvOJDcruayagGA6wu9hRrTUpOtjrQG4ZoqUGe
DSBZk/VDAE2TO4BcXhlyyBdY0Wt5rMW1jDO71bRCaHIQpOMPhDs3ad1uxPkbsiCS
GfNSrUe81gN89LYWt+2jy3hHOQuPjHqvedqnmqOcpdi8zuQFYQSGmq83ZK2hnnWa
3pDmWKgpEOAtQ1H5LBxnhF44O6SlWAFoGe2rBf2v6DqsNHi/iWy+Ry+OVRQHRzmi
QMmH7BdsjXpnuRzai9qNHyWUf70SL5mKGUN7yIWl4bQ8CzBpStQRzOgJLSvz6V5E
Im/20KcUMklXf58Fqc8+FJCzHsAAhT091qqILQTyDZOPYl36Kh2j4M2JIHKT4CcE
XJoZTEMhuaYlzVqKRq4RfN6XrObbfaLp9NRBlr94HqaU1oyf5vBL8hGPDaI96bI+
7cWxpXh0LVHezCFLMY57Qal9svMLtpTgiAwEAZSpjePJXn5TB+8LOMxlMTilPDzY
lndzL0PLCB0dXOc0BXFn6CajeYnbgF5mZdAwteDsoyFOZyeS9YvS1OEQgIsMAoIV
0+cnrHzgG0YvMcu8WX/xgAEZeMdx00f0xcRk3RJ5AnX4r4NW+rJDpq137uerZCIQ
cRPAdo95xl14Yn4FMc4S5FcWxDJUMCZKJFPPNCC58RNeAZA0eFSsEzcsAakOR52W
OHD0XNQaIc0qOeDJOJIkNA+VIfQsi4mpqETgmemZNJ3lnJo33Rfl4jooxQPoYXY0
xylNr7OXfHH96q83v5ugcR8T90gHi2QfrGBrkVcCLjPjYEhk8O4xTXOIANd/Ca6t
Uzp7KczvV/buNWbSmR9KwkH281Ernv7BYAmKOjotw4dFvCovnWHQqvIOxNbIa0H2
hGQj/i4o6Y43Co7Ln4+v8ud9lvWsg3TiSEcC7EYc0O/NWDJi81byIxXw1UrS5oKQ
g8AZs3LnzttVganSyYwrX0Fnk57L249O2lES4w7F7kvoABNihzcjQ5GYCZE6HfJv
Zvjxu8hZPRfMkuDiZh4EUkkxmZqaUJzkhzD3RUzWQ0sJWeMxTjfW/2FZTA9adktM
rgxCXT/8ShhRU5rxWuB+4CC2s2PxeygCfdixyKNeiYTL3+kA9dsQLqoKNxX7wWgJ
0X4RZJ3LqBNSN/NmgcvPOa8rxilpaCCSecnErw/MtYzmNhQM78LUkYXWd5eV64fc
dngvvIgiQk4e0fhzsCPyFIJkYa1UKKCI0Ye4342KLcTuB9n4hz8MV5uMtnxeEq3K
5aXgGRRNkcKjmd7FnQ2hy0U8K2zj9SHvCFHEpeln7IUPKKoJc307O2yM8wbYcWpY
K7gw3O6I3Y0d2dKHqKqpR40Yalysn0seTdRga9C/9jnkVbnxBH8ne/VKeK6aII+B
xse/Pb2N/Je6GKqpdsnXa1jRs17+iMqh5JuiJVGYmmOX4JekIs6UTf5zV/4p6Nse
iMjM7HrRnISRv8w4nLQCXxYyukelUfN0bJbdZjX1JELdlkS5awNcO0XWOTxKfaoV
Mw+2cVlPz8IdsMHJjviY9eeESmobCbgj5fsbShQMfuTvvmY1PgeEcmjgn1DjWfrq
0QebnnbQEY63mtQyjyteej+4RMrzjZoZFBfY1DFcnrV1oxQ4LtA9Y2IM8BnrTON3
Q784F3cEQzqEy8/qKAyJfl+wfK+6q1wM/v/DjJySw5tu/NPgYrHrYdn5pP+/r69h
o3mcFqgKjBHK8qhV+t/qG2o7TkL25fIwhilQa33jHCCTgz0Q7Wf43bfvPQflRYqz
u1zjGOHK/ghmnATFQkf04y3KycveGYFjDZ8+rmVlFqGPRBgwc0s+ifqpAV7cW8jA
/NTB+Am8LuJ8rT/QkrjXwTLextXtSIig6PggpN8tYjeenY1Z7QunGHvMjYGPHcm/
S/lkR3uunF/Xj7aMTm/p+Wtom8DjCCTZDEIN2vmuzsKNHp7899I3DNutiCxXv4b8
0cJFrlvZuYZ6z32w9WA6EZB1pJ5e6ra+ZInzKJYLgc/OWbo93u3w2X+sn3FnfoQO
8T6NbGwdm7fNBNhBFO7saozXWI+WhyGjTvsJaeRBZmA2FbM7wNX0G9dTyF6ns96b
rVZs+hZjNmiBTDWO1QPJPzhbQ4fqNymLtgHDG2/VP839qOj6NHqApJC0OSH8YOnk
e8B4b8/iFrpdBtHqbRq9sn9/l0RxrNLVvUZAexG4D/QxVRfPAs6HO23Qqahb4/16
WNqFZLYuDJ/++1MXDT1JaLuVWkTqi3Lh/1NCFEt5Rf5fbgJWhj54Drw5z2H/NdnC
hhmC0u6CazXOgD0TnOI2IO5ERdFq06hssjKjrNmNb9TNr9FL62Bzf+vhHYyCF704
KvenXtuBe9dE5Vc9IHxD5nWX5RUiTvgiSAygaLVJdbXX4WjwyvLf7ErMXdudunNN
vw2RNEIx0GJeaQDgZwY4nmZt4xKfsiabVp+kjsvGLwEDdQtj+aS31Pagzxen0I5n
2IBEGNjXEc+pTIVJgiVGEueiLpcnTPo+YVkVA+nIUY0FMPk+pekpUL2ixAczsRdW
Hn/GgIS93kvAsSMkADhZe47xmG0/Kz/nRCW9vGz2551Xh8EkXig5RNL+F+5rHs5a
te95atJ9aqmrxYeClx05ncYpkkueMtXk7aE1qDF0rJtKaS1+nv4IhCAocS+dRo1q
7PoArdZ/rlDNjw8i1KsqaFES0kC6o7kUwhMMD1txbITvemclx6w0BoQU4A3cf6If
QoTPBAAany9RrtZ+niebE7RQEZRJJLuFLEYeIxgBN7/9ovguZDDLadTTTvWESzs4
RsjEy2GvEAvYGN83QXNp99FEs+dfr5jshdjlo454LuCCQviCzntp67trKQx9kMqU
FKQ00zOP/eNIOS6Ojh581INHGARMyfgHdblhLgMWoiXCWNzP4qOiHCa/D+yEiTjF
G1DkoGDuxo76SIuq0vAK6RjWYkcCLt8/TlMCSyPfcPKGJNbgRJesNp6JI8BsNc5N
aItbZNmQo9rbTuAAFKibEQ8DACZcaJEbyNXZ6lx97/uWNw8mPIB7vp2el+al8/YI
xvPNSsRUcbJ2Kz8bD2sfpE7tzFRvXs0o8zt0oyKjUrPNAHntRcz19WTA8bua8Ez6
0SREk9uaGIfl7PEyID/gjmdVB4OIUD0H6BjMb99yBFStFDzpeM3qVd6ivYVw9k1u
Z2g0rgijagrPtN5QJsikjUlgQQE00vOd0HSv6RtK2YrHhBrBhFlSZuXr32jzFw1A
nZl9d95hx9EVm0em5GE/D14jwFwEUzQdXiFwJQt+V2UMWvdfW/kQQBKfRGOaC3GU
jdMNGv9peg5rRw9yRzyTa8GS67Q/ggnU/l/y7l5ecapFVhVH5IdPNHVAz+roc6pP
Y9iIxeWRQijEBfSumC9iN7LHmkdjmUOCtClW7uC9H+BXDyNrLliRtryb+F/wGTzH
ZgVv4l3pdAu2WSP9x+5lmAXAvKKhuKXLcX9mVIP8Mk1n2dn3HxCzC7TrHuZ2c0dd
Q+7yPz2yxn3u7a6HWyiiSymTyWCIesQ03OsOzug4CwHK6hD3kWiklA+fOexr0jZ6
4xlauYpSVv4UjltClvrXgeuQBCFjj/PrcwEE0yfAyqkMh7ykROpgbU2H5CFaqcXB
BDJApcay3VpegIMkBQXnYkGcz6a1fnzTMJP85q8SkMBwlqLqo+X7uRrt4VXwVt+/
oizl/NAio0geu4IVywPYUdVkWdlaxbNgU/T3dWUyI8RmwqPU82dulcj1zCLUtw6d
EQaiT4c9xKtXXNhHN5Hty6f1Hj4evTfWnaGb/PxZD0og9x+ns95RDMEm381kHoQP
nIURAEcyRU66jVVoJn3jLVTFLwotJqzZ17WnfRad/Gy0M0yLEyeXtywdVxo9I6D0
siO9XwE0YYWCE6QYwzJpwyS/97X4xFGFGIvswDQ8u927DqVRUS51jJeWD+dZrccw
/navSCS38Ho+O8WEWeAEPjCAQmC1ukMtkRIdUMwMlGcu2NewdjjVKO+e22D7oJe1
VCB+AYRwZxoQM3D20e5DFSYdLR3YF6SiutVUlbwntdt0BGIIIdgjBAVXb+j2qwn+
WTfKKzbJW0v4rrx6PxvGEYMYEBbUFICwgylhBYQCziEwrIQsrRoclWI8Sr731urK
mxDC2nMVbECOdqw/roZ+XhoYqICu8A0+e9tYa8R+irmGIdoIR/eKhBOxlwwN8dDS
mY2A8mSsyj/or/LVyqPDGQ51FHeuLKWrXMFKLyP6DTRumrmFBhMD8lTRrpa5/2TG
eA1vm5lhyLYBWLo1GYlkhQq4o+5M4vRuu6KlLZEk9gsDOUoqEczGqvNMQpFX8aME
qvu8U/nEl1F2YdAurb6whALjDetXur7qfYwS8NkHfVTXsVlu8rKr8dWnBYjREt3s
DN9Be1UE3glkzolUt7MIzwpnJIX1XTXvUBwovsk7QI4lSzBtUZ2PgrH6Yx2kz0Z9
lGzxBWFSLtCzgjkV3tlB/DqodIGOQ939IknemsOmN+Jr5HJdbN33ecydOFQ+3Gq9
ZqnPQ8Pah8l/IyS0UaCmu3AIGiswd0W8MAbrHDtQFIsxWIMLr81TFdsKu31C0q0S
PohxAuuASyymxc3C8KcfQOgepqN1bgVIT/WjocPooagi6dypXGjBz+3KW6aMR1Co
xu8iM2GFbSrs6FHG24O5ebFyVbCNGaLg9nMEYophlaKl8JTuprKcRU7f7vR35Fbk
hICoGRZYw+63FH0jus/FlNZqFlqFxADxL3giqfJtyMZNhwGfTcaOdlNVonjI764h
DXoT6HO0zULJUfFzXQHQ6+RICft7EUBOBVOIdckN9PKFi9An3uNKOBduyCanVABL
0orOxnZp+9uT+LbrBCBzNcw928mQsnUrFpDNp1yYULrldgl5ZIXJbuDKlwngVUiS
ebc2ELowIoX3JvDrguGoWPRrTBdX5AxbsRU0Lz6LQ1Tc0s4s9piG7v+vbVFQ/UEL
Lbhnes68Wpa1ZvHV9MALskaZLA6S/Jles6YW60Ke0BYWF5VZXLFXFkoddI5UcgQF
8DMwimQCgZiLwq47D/WD7fvFzR2A/d29zmvfJrOEv2ccQVC7j1MPTEoK4yFWSAmf
ll6/Z1bfmNnopo4pk+wbodaztNjhLQg07Ed2xLaALt2/xmFOY3DNscCTuN/Zc8FF
DV/zY6ikjaR05Tct4yYvI7kXFHf5LsBWqGcE5KRBCeFDPsX9c5XEWU1KYyastMfN
Vo1ZZ+F7dSUmTMbzMbZoUEIiix/Sc5A16TzmfV734a7NkLOuE7tuQHhlBQULt4Sq
jaxcOfMw6cv6I20FYmIWW39rOUUlF/sMc0PDvsL9v7yGEjh9eeFuLWxmEBlG7TEb
XdDYMENSabCIJBNsWg1eRGgDA+FWvBCVVnUnfLkcof33e0Y3eLj8D8f0x6bfAPQe
hTWtu4bxptQ7ua6wYJknysVS9x4bVSOl/vnbeHqfTezPQrL6CfBaAD3HX0gFxvMZ
KLMnFTe+wXtgX18f32tUSaLMnXyGZ+WLHol9bH31y8AWB6EL+oOeDcS7WOybgzYs
F0TgBpztufbsn1CiICOm9S5QCH9vv4GIggTK9vb8Zu2w6VP3BaHdDeeNNCc2dp2f
0xnHchomFxvbR/kRlA5Cg4wq8kK9WZNmACbdAek5pDy8i0WYmx46sMahjXRXnTU5
+gOOv5UkcaYhOKmP6HGt3xIIcsAifmgxHYkvsehFaRTvDMLKNfKHQDazVKuNXk/E
hoWj+Wk5LwVOvEgNljTC2Uz/wpo8xW+Fmp7hyKX4t5m2PHOKwDWDnjKmLED73Vf4
RdKtAIbkLJP90i68Jsb52eMRW2IU/ne/g7F0swXn+qo3eyR6QKYw9I4Q8t0hjxiI
IraCY4Qa3BBXINCBY+i+XFmjNZdaY3l0+F5ujQpVWfFZ7RiWiGt0k7hvTsAUvX2c
SZtwEYTkNRKW1SRlqvLhFGfmhoUQk7Qai3h6bwLFV5U=
//pragma protect end_data_block
//pragma protect digest_block
gpzroK1hTR5sY30DqW4rHFPJdYY=
//pragma protect end_digest_block
//pragma protect end_protected
`endprotect
