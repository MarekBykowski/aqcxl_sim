`protected
TWBg.?-)XDFg8-aQbW<bM&Y]>ZL[_<e&\?Q??.GRZeJ):/5f00BK/)/eR1]:@+_+
WH+&5DH1a1F(A(\PfD<7&/^_Qf56^bV)GZ/3PU?E/,34E;.ZgJ;e=QUa0c<#,VYJ
:9?8^f6E?^C\_8WC#ERBZTSg5f0Z:L.E<TF0g=ET[Y=2942aJ,DXcABAVU^ILb)6
dT5<O[F.UB;9dg>7SEFE^B0A)@gA8cCT-]N]OVXP:C2UFIeL5N&aFZA8>KS;cIbP
9T^^1K?bf0d;O2/AF92U>VHX/;(N6STf]RbIO5YFXL8&C[e(5O2B;B)fK<7OS-Ze
,d@X-=^Y.A2;*$
`endprotected

